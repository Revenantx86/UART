VERSION 5.8 ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;
UNITS
    DATABASE MICRONS 1000 ;
END UNITS

VIA via2_3_2000_480_1_6_320_320
  VIARULE M1M2_PR ;
  CUTSIZE 0.15 0.15 ;
  LAYERS met1 via met2 ;
  CUTSPACING 0.17 0.17 ;
  ENCLOSURE 0.085 0.165 0.055 0.085 ;
  ROWCOL 1 6 ;
END via2_3_2000_480_1_6_320_320

VIA via3_4_2000_480_1_5_400_400
  VIARULE M2M3_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met2 via2 met3 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.04 0.085 0.065 0.065 ;
  ROWCOL 1 5 ;
END via3_4_2000_480_1_5_400_400

VIA via4_5_2000_480_1_5_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.06 0.1 0.065 ;
  ROWCOL 1 5 ;
END via4_5_2000_480_1_5_400_400

VIA via4_5_2000_2000_5_5_400_400
  VIARULE M3M4_PR ;
  CUTSIZE 0.2 0.2 ;
  LAYERS met3 via3 met4 ;
  CUTSPACING 0.2 0.2 ;
  ENCLOSURE 0.09 0.1 0.1 0.065 ;
  ROWCOL 5 5 ;
END via4_5_2000_2000_5_5_400_400

MACRO fifo
  FOREIGN fifo 0 0 ;
  CLASS BLOCK ;
  SIZE 128.98 BY 247.36 ;
  PIN VSS
    USE GROUND ;
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT  1.38 236.4 124.98 236.88 ;
        RECT  1.38 230.96 124.98 231.44 ;
        RECT  1.38 225.52 124.98 226 ;
        RECT  1.38 220.08 124.98 220.56 ;
        RECT  1.38 214.64 124.98 215.12 ;
        RECT  1.38 209.2 124.98 209.68 ;
        RECT  1.38 203.76 124.98 204.24 ;
        RECT  1.38 198.32 124.98 198.8 ;
        RECT  1.38 192.88 124.98 193.36 ;
        RECT  1.38 187.44 124.98 187.92 ;
        RECT  1.38 182 124.98 182.48 ;
        RECT  1.38 176.56 124.98 177.04 ;
        RECT  1.38 171.12 124.98 171.6 ;
        RECT  1.38 165.68 124.98 166.16 ;
        RECT  1.38 160.24 124.98 160.72 ;
        RECT  1.38 154.8 124.98 155.28 ;
        RECT  1.38 149.36 124.98 149.84 ;
        RECT  1.38 143.92 124.98 144.4 ;
        RECT  1.38 138.48 124.98 138.96 ;
        RECT  1.38 133.04 124.98 133.52 ;
        RECT  1.38 127.6 124.98 128.08 ;
        RECT  1.38 122.16 124.98 122.64 ;
        RECT  1.38 116.72 124.98 117.2 ;
        RECT  1.38 111.28 124.98 111.76 ;
        RECT  1.38 105.84 124.98 106.32 ;
        RECT  1.38 100.4 124.98 100.88 ;
        RECT  1.38 94.96 124.98 95.44 ;
        RECT  1.38 89.52 124.98 90 ;
        RECT  1.38 84.08 124.98 84.56 ;
        RECT  1.38 78.64 124.98 79.12 ;
        RECT  1.38 73.2 124.98 73.68 ;
        RECT  1.38 67.76 124.98 68.24 ;
        RECT  1.38 62.32 124.98 62.8 ;
        RECT  1.38 56.88 124.98 57.36 ;
        RECT  1.38 51.44 124.98 51.92 ;
        RECT  1.38 46 124.98 46.48 ;
        RECT  1.38 40.56 124.98 41.04 ;
        RECT  1.38 35.12 124.98 35.6 ;
        RECT  1.38 29.68 124.98 30.16 ;
        RECT  1.38 24.24 124.98 24.72 ;
        RECT  1.38 18.8 124.98 19.28 ;
        RECT  1.38 13.36 124.98 13.84 ;
        RECT  1.38 7.92 124.98 8.4 ;
        RECT  1.38 2.48 124.98 2.96 ;
      LAYER met4 ;
        RECT  122.98 -1.28 124.98 243.36 ;
      LAYER met3 ;
        RECT  -2.62 241.36 124.98 243.36 ;
        RECT  -2.62 -1.28 124.98 0.72 ;
      LAYER met4 ;
        RECT  -2.62 -1.28 -0.62 243.36 ;
      VIA 123.98 242.36 via4_5_2000_2000_5_5_400_400 ;
      VIA 123.98 -0.28 via4_5_2000_2000_5_5_400_400 ;
      VIA -1.62 242.36 via4_5_2000_2000_5_5_400_400 ;
      VIA -1.62 -0.28 via4_5_2000_2000_5_5_400_400 ;
      LAYER met3 ;
        RECT  122.99 236.475 124.97 236.805 ;
      VIA 123.98 236.64 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 236.64 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 236.64 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 231.035 124.97 231.365 ;
      VIA 123.98 231.2 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 231.2 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 231.2 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 225.595 124.97 225.925 ;
      VIA 123.98 225.76 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 225.76 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 225.76 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 220.155 124.97 220.485 ;
      VIA 123.98 220.32 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 220.32 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 220.32 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 214.715 124.97 215.045 ;
      VIA 123.98 214.88 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 214.88 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 214.88 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 209.275 124.97 209.605 ;
      VIA 123.98 209.44 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 209.44 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 209.44 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 203.835 124.97 204.165 ;
      VIA 123.98 204 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 204 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 204 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 198.395 124.97 198.725 ;
      VIA 123.98 198.56 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 198.56 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 198.56 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 192.955 124.97 193.285 ;
      VIA 123.98 193.12 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 193.12 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 193.12 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 187.515 124.97 187.845 ;
      VIA 123.98 187.68 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 187.68 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 187.68 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 182.075 124.97 182.405 ;
      VIA 123.98 182.24 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 182.24 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 182.24 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 176.635 124.97 176.965 ;
      VIA 123.98 176.8 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 176.8 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 176.8 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 171.195 124.97 171.525 ;
      VIA 123.98 171.36 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 171.36 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 171.36 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 165.755 124.97 166.085 ;
      VIA 123.98 165.92 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 165.92 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 165.92 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 160.315 124.97 160.645 ;
      VIA 123.98 160.48 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 160.48 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 160.48 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 154.875 124.97 155.205 ;
      VIA 123.98 155.04 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 155.04 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 155.04 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 149.435 124.97 149.765 ;
      VIA 123.98 149.6 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 149.6 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 149.6 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 143.995 124.97 144.325 ;
      VIA 123.98 144.16 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 144.16 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 144.16 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 138.555 124.97 138.885 ;
      VIA 123.98 138.72 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 138.72 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 138.72 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 133.115 124.97 133.445 ;
      VIA 123.98 133.28 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 133.28 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 133.28 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 127.675 124.97 128.005 ;
      VIA 123.98 127.84 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 127.84 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 127.84 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 122.235 124.97 122.565 ;
      VIA 123.98 122.4 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 122.4 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 122.4 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 116.795 124.97 117.125 ;
      VIA 123.98 116.96 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 116.96 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 116.96 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 111.355 124.97 111.685 ;
      VIA 123.98 111.52 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 111.52 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 111.52 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 105.915 124.97 106.245 ;
      VIA 123.98 106.08 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 106.08 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 106.08 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 100.475 124.97 100.805 ;
      VIA 123.98 100.64 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 100.64 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 100.64 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 95.035 124.97 95.365 ;
      VIA 123.98 95.2 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 95.2 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 95.2 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 89.595 124.97 89.925 ;
      VIA 123.98 89.76 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 89.76 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 89.76 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 84.155 124.97 84.485 ;
      VIA 123.98 84.32 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 84.32 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 84.32 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 78.715 124.97 79.045 ;
      VIA 123.98 78.88 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 78.88 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 78.88 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 73.275 124.97 73.605 ;
      VIA 123.98 73.44 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 73.44 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 73.44 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 67.835 124.97 68.165 ;
      VIA 123.98 68 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 68 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 68 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 62.395 124.97 62.725 ;
      VIA 123.98 62.56 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 62.56 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 62.56 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 56.955 124.97 57.285 ;
      VIA 123.98 57.12 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 57.12 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 57.12 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 51.515 124.97 51.845 ;
      VIA 123.98 51.68 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 51.68 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 51.68 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 46.075 124.97 46.405 ;
      VIA 123.98 46.24 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 46.24 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 46.24 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 40.635 124.97 40.965 ;
      VIA 123.98 40.8 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 40.8 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 40.8 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 35.195 124.97 35.525 ;
      VIA 123.98 35.36 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 35.36 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 35.36 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 29.755 124.97 30.085 ;
      VIA 123.98 29.92 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 29.92 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 29.92 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 24.315 124.97 24.645 ;
      VIA 123.98 24.48 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 24.48 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 24.48 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 18.875 124.97 19.205 ;
      VIA 123.98 19.04 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 19.04 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 19.04 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 13.435 124.97 13.765 ;
      VIA 123.98 13.6 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 13.6 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 13.6 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 7.995 124.97 8.325 ;
      VIA 123.98 8.16 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 8.16 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 8.16 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  122.99 2.555 124.97 2.885 ;
      VIA 123.98 2.72 via4_5_2000_480_1_5_400_400 ;
      VIA 123.98 2.72 via3_4_2000_480_1_5_400_400 ;
      VIA 123.98 2.72 via2_3_2000_480_1_6_320_320 ;
    END
  END VSS
  PIN VDD
    USE POWER ;
    DIRECTION INOUT ;
    PORT
      LAYER met1 ;
        RECT  -6.62 239.12 128.98 239.6 ;
        RECT  -6.62 233.68 128.98 234.16 ;
        RECT  -6.62 228.24 128.98 228.72 ;
        RECT  -6.62 222.8 128.98 223.28 ;
        RECT  -6.62 217.36 128.98 217.84 ;
        RECT  -6.62 211.92 128.98 212.4 ;
        RECT  -6.62 206.48 128.98 206.96 ;
        RECT  -6.62 201.04 128.98 201.52 ;
        RECT  -6.62 195.6 128.98 196.08 ;
        RECT  -6.62 190.16 128.98 190.64 ;
        RECT  -6.62 184.72 128.98 185.2 ;
        RECT  -6.62 179.28 128.98 179.76 ;
        RECT  -6.62 173.84 128.98 174.32 ;
        RECT  -6.62 168.4 128.98 168.88 ;
        RECT  -6.62 162.96 128.98 163.44 ;
        RECT  -6.62 157.52 128.98 158 ;
        RECT  -6.62 152.08 128.98 152.56 ;
        RECT  -6.62 146.64 128.98 147.12 ;
        RECT  -6.62 141.2 128.98 141.68 ;
        RECT  -6.62 135.76 128.98 136.24 ;
        RECT  -6.62 130.32 128.98 130.8 ;
        RECT  -6.62 124.88 128.98 125.36 ;
        RECT  -6.62 119.44 128.98 119.92 ;
        RECT  -6.62 114 128.98 114.48 ;
        RECT  -6.62 108.56 128.98 109.04 ;
        RECT  -6.62 103.12 128.98 103.6 ;
        RECT  -6.62 97.68 128.98 98.16 ;
        RECT  -6.62 92.24 128.98 92.72 ;
        RECT  -6.62 86.8 128.98 87.28 ;
        RECT  -6.62 81.36 128.98 81.84 ;
        RECT  -6.62 75.92 128.98 76.4 ;
        RECT  -6.62 70.48 128.98 70.96 ;
        RECT  -6.62 65.04 128.98 65.52 ;
        RECT  -6.62 59.6 128.98 60.08 ;
        RECT  -6.62 54.16 128.98 54.64 ;
        RECT  -6.62 48.72 128.98 49.2 ;
        RECT  -6.62 43.28 128.98 43.76 ;
        RECT  -6.62 37.84 128.98 38.32 ;
        RECT  -6.62 32.4 128.98 32.88 ;
        RECT  -6.62 26.96 128.98 27.44 ;
        RECT  -6.62 21.52 128.98 22 ;
        RECT  -6.62 16.08 128.98 16.56 ;
        RECT  -6.62 10.64 128.98 11.12 ;
        RECT  -6.62 5.2 128.98 5.68 ;
      LAYER met4 ;
        RECT  126.98 -5.28 128.98 247.36 ;
      LAYER met3 ;
        RECT  -6.62 245.36 128.98 247.36 ;
        RECT  -6.62 -5.28 128.98 -3.28 ;
      LAYER met4 ;
        RECT  -6.62 -5.28 -4.62 247.36 ;
      VIA 127.98 246.36 via4_5_2000_2000_5_5_400_400 ;
      VIA 127.98 -4.28 via4_5_2000_2000_5_5_400_400 ;
      VIA -5.62 246.36 via4_5_2000_2000_5_5_400_400 ;
      VIA -5.62 -4.28 via4_5_2000_2000_5_5_400_400 ;
      LAYER met3 ;
        RECT  126.99 239.195 128.97 239.525 ;
      VIA 127.98 239.36 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 239.36 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 239.36 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 233.755 128.97 234.085 ;
      VIA 127.98 233.92 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 233.92 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 233.92 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 228.315 128.97 228.645 ;
      VIA 127.98 228.48 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 228.48 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 228.48 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 222.875 128.97 223.205 ;
      VIA 127.98 223.04 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 223.04 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 223.04 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 217.435 128.97 217.765 ;
      VIA 127.98 217.6 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 217.6 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 217.6 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 211.995 128.97 212.325 ;
      VIA 127.98 212.16 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 212.16 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 212.16 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 206.555 128.97 206.885 ;
      VIA 127.98 206.72 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 206.72 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 206.72 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 201.115 128.97 201.445 ;
      VIA 127.98 201.28 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 201.28 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 201.28 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 195.675 128.97 196.005 ;
      VIA 127.98 195.84 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 195.84 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 195.84 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 190.235 128.97 190.565 ;
      VIA 127.98 190.4 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 190.4 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 190.4 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 184.795 128.97 185.125 ;
      VIA 127.98 184.96 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 184.96 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 184.96 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 179.355 128.97 179.685 ;
      VIA 127.98 179.52 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 179.52 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 179.52 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 173.915 128.97 174.245 ;
      VIA 127.98 174.08 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 174.08 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 174.08 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 168.475 128.97 168.805 ;
      VIA 127.98 168.64 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 168.64 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 168.64 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 163.035 128.97 163.365 ;
      VIA 127.98 163.2 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 163.2 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 163.2 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 157.595 128.97 157.925 ;
      VIA 127.98 157.76 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 157.76 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 157.76 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 152.155 128.97 152.485 ;
      VIA 127.98 152.32 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 152.32 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 152.32 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 146.715 128.97 147.045 ;
      VIA 127.98 146.88 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 146.88 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 146.88 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 141.275 128.97 141.605 ;
      VIA 127.98 141.44 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 141.44 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 141.44 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 135.835 128.97 136.165 ;
      VIA 127.98 136 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 136 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 136 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 130.395 128.97 130.725 ;
      VIA 127.98 130.56 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 130.56 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 130.56 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 124.955 128.97 125.285 ;
      VIA 127.98 125.12 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 125.12 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 125.12 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 119.515 128.97 119.845 ;
      VIA 127.98 119.68 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 119.68 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 119.68 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 114.075 128.97 114.405 ;
      VIA 127.98 114.24 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 114.24 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 114.24 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 108.635 128.97 108.965 ;
      VIA 127.98 108.8 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 108.8 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 108.8 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 103.195 128.97 103.525 ;
      VIA 127.98 103.36 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 103.36 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 103.36 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 97.755 128.97 98.085 ;
      VIA 127.98 97.92 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 97.92 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 97.92 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 92.315 128.97 92.645 ;
      VIA 127.98 92.48 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 92.48 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 92.48 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 86.875 128.97 87.205 ;
      VIA 127.98 87.04 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 87.04 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 87.04 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 81.435 128.97 81.765 ;
      VIA 127.98 81.6 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 81.6 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 81.6 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 75.995 128.97 76.325 ;
      VIA 127.98 76.16 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 76.16 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 76.16 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 70.555 128.97 70.885 ;
      VIA 127.98 70.72 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 70.72 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 70.72 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 65.115 128.97 65.445 ;
      VIA 127.98 65.28 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 65.28 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 65.28 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 59.675 128.97 60.005 ;
      VIA 127.98 59.84 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 59.84 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 59.84 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 54.235 128.97 54.565 ;
      VIA 127.98 54.4 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 54.4 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 54.4 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 48.795 128.97 49.125 ;
      VIA 127.98 48.96 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 48.96 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 48.96 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 43.355 128.97 43.685 ;
      VIA 127.98 43.52 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 43.52 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 43.52 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 37.915 128.97 38.245 ;
      VIA 127.98 38.08 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 38.08 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 38.08 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 32.475 128.97 32.805 ;
      VIA 127.98 32.64 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 32.64 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 32.64 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 27.035 128.97 27.365 ;
      VIA 127.98 27.2 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 27.2 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 27.2 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 21.595 128.97 21.925 ;
      VIA 127.98 21.76 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 21.76 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 21.76 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 16.155 128.97 16.485 ;
      VIA 127.98 16.32 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 16.32 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 16.32 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 10.715 128.97 11.045 ;
      VIA 127.98 10.88 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 10.88 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 10.88 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  126.99 5.275 128.97 5.605 ;
      VIA 127.98 5.44 via4_5_2000_480_1_5_400_400 ;
      VIA 127.98 5.44 via3_4_2000_480_1_5_400_400 ;
      VIA 127.98 5.44 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 239.195 -4.63 239.525 ;
      VIA -5.62 239.36 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 239.36 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 239.36 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 233.755 -4.63 234.085 ;
      VIA -5.62 233.92 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 233.92 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 233.92 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 228.315 -4.63 228.645 ;
      VIA -5.62 228.48 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 228.48 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 228.48 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 222.875 -4.63 223.205 ;
      VIA -5.62 223.04 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 223.04 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 223.04 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 217.435 -4.63 217.765 ;
      VIA -5.62 217.6 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 217.6 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 217.6 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 211.995 -4.63 212.325 ;
      VIA -5.62 212.16 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 212.16 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 212.16 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 206.555 -4.63 206.885 ;
      VIA -5.62 206.72 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 206.72 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 206.72 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 201.115 -4.63 201.445 ;
      VIA -5.62 201.28 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 201.28 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 201.28 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 195.675 -4.63 196.005 ;
      VIA -5.62 195.84 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 195.84 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 195.84 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 190.235 -4.63 190.565 ;
      VIA -5.62 190.4 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 190.4 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 190.4 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 184.795 -4.63 185.125 ;
      VIA -5.62 184.96 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 184.96 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 184.96 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 179.355 -4.63 179.685 ;
      VIA -5.62 179.52 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 179.52 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 179.52 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 173.915 -4.63 174.245 ;
      VIA -5.62 174.08 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 174.08 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 174.08 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 168.475 -4.63 168.805 ;
      VIA -5.62 168.64 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 168.64 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 168.64 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 163.035 -4.63 163.365 ;
      VIA -5.62 163.2 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 163.2 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 163.2 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 157.595 -4.63 157.925 ;
      VIA -5.62 157.76 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 157.76 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 157.76 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 152.155 -4.63 152.485 ;
      VIA -5.62 152.32 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 152.32 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 152.32 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 146.715 -4.63 147.045 ;
      VIA -5.62 146.88 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 146.88 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 146.88 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 141.275 -4.63 141.605 ;
      VIA -5.62 141.44 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 141.44 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 141.44 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 135.835 -4.63 136.165 ;
      VIA -5.62 136 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 136 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 136 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 130.395 -4.63 130.725 ;
      VIA -5.62 130.56 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 130.56 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 130.56 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 124.955 -4.63 125.285 ;
      VIA -5.62 125.12 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 125.12 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 125.12 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 119.515 -4.63 119.845 ;
      VIA -5.62 119.68 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 119.68 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 119.68 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 114.075 -4.63 114.405 ;
      VIA -5.62 114.24 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 114.24 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 114.24 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 108.635 -4.63 108.965 ;
      VIA -5.62 108.8 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 108.8 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 108.8 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 103.195 -4.63 103.525 ;
      VIA -5.62 103.36 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 103.36 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 103.36 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 97.755 -4.63 98.085 ;
      VIA -5.62 97.92 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 97.92 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 97.92 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 92.315 -4.63 92.645 ;
      VIA -5.62 92.48 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 92.48 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 92.48 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 86.875 -4.63 87.205 ;
      VIA -5.62 87.04 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 87.04 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 87.04 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 81.435 -4.63 81.765 ;
      VIA -5.62 81.6 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 81.6 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 81.6 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 75.995 -4.63 76.325 ;
      VIA -5.62 76.16 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 76.16 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 76.16 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 70.555 -4.63 70.885 ;
      VIA -5.62 70.72 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 70.72 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 70.72 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 65.115 -4.63 65.445 ;
      VIA -5.62 65.28 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 65.28 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 65.28 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 59.675 -4.63 60.005 ;
      VIA -5.62 59.84 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 59.84 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 59.84 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 54.235 -4.63 54.565 ;
      VIA -5.62 54.4 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 54.4 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 54.4 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 48.795 -4.63 49.125 ;
      VIA -5.62 48.96 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 48.96 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 48.96 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 43.355 -4.63 43.685 ;
      VIA -5.62 43.52 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 43.52 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 43.52 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 37.915 -4.63 38.245 ;
      VIA -5.62 38.08 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 38.08 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 38.08 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 32.475 -4.63 32.805 ;
      VIA -5.62 32.64 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 32.64 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 32.64 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 27.035 -4.63 27.365 ;
      VIA -5.62 27.2 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 27.2 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 27.2 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 21.595 -4.63 21.925 ;
      VIA -5.62 21.76 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 21.76 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 21.76 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 16.155 -4.63 16.485 ;
      VIA -5.62 16.32 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 16.32 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 16.32 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 10.715 -4.63 11.045 ;
      VIA -5.62 10.88 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 10.88 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 10.88 via2_3_2000_480_1_6_320_320 ;
      LAYER met3 ;
        RECT  -6.61 5.275 -4.63 5.605 ;
      VIA -5.62 5.44 via4_5_2000_480_1_5_400_400 ;
      VIA -5.62 5.44 via3_4_2000_480_1_5_400_400 ;
      VIA -5.62 5.44 via2_3_2000_480_1_6_320_320 ;
    END
  END VDD
  PIN clk
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 232.75 0.8 233.05 ;
    END
  END clk
  PIN data_in[0]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 213.71 0.8 214.01 ;
    END
  END data_in[0]
  PIN data_in[1]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  93.08 241.95 93.22 242.435 ;
    END
  END data_in[1]
  PIN data_in[2]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 231.39 0.8 231.69 ;
    END
  END data_in[2]
  PIN data_in[3]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  121.415 8.35 122.215 8.65 ;
    END
  END data_in[3]
  PIN data_in[4]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  121.415 26.03 122.215 26.33 ;
    END
  END data_in[4]
  PIN data_in[5]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  106.88 241.95 107.02 242.435 ;
    END
  END data_in[5]
  PIN data_in[6]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  121.415 9.71 122.215 10.01 ;
    END
  END data_in[6]
  PIN data_in[7]
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  110.56 241.95 110.7 242.435 ;
    END
  END data_in[7]
  PIN data_out[0]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 129.39 0.8 129.69 ;
    END
  END data_out[0]
  PIN data_out[1]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 144.35 0.8 144.65 ;
    END
  END data_out[1]
  PIN data_out[2]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 141.63 0.8 141.93 ;
    END
  END data_out[2]
  PIN data_out[3]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 113.07 0.8 113.37 ;
    END
  END data_out[3]
  PIN data_out[4]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 126.67 0.8 126.97 ;
    END
  END data_out[4]
  PIN data_out[5]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 114.43 0.8 114.73 ;
    END
  END data_out[5]
  PIN data_out[6]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 140.27 0.8 140.57 ;
    END
  END data_out[6]
  PIN data_out[7]
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 142.99 0.8 143.29 ;
    END
  END data_out[7]
  PIN empty
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  2.92 241.95 3.06 242.435 ;
    END
  END empty
  PIN full
    DIRECTION OUTPUT ;
    USE SIGNAL ;
    PORT
      LAYER met2 ;
        RECT  3.84 241.95 3.98 242.435 ;
    END
  END full
  PIN rd_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 110.35 0.8 110.65 ;
    END
  END rd_en
  PIN rst
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  0 108.99 0.8 109.29 ;
    END
  END rst
  PIN wr_en
    DIRECTION INPUT ;
    USE SIGNAL ;
    PORT
      LAYER met3 ;
        RECT  121.415 74.99 122.215 75.29 ;
    END
  END wr_en
  OBS
    LAYER nwell ;
     RECT  1.19 4.025 121.17 6.855 ;
     RECT  1.19 9.465 121.17 12.295 ;
     RECT  1.19 14.905 121.17 17.735 ;
     RECT  1.19 20.345 121.17 23.175 ;
     RECT  1.19 25.785 121.17 28.615 ;
     RECT  1.19 31.225 121.17 34.055 ;
     RECT  1.19 36.665 121.17 39.495 ;
     RECT  1.19 42.105 121.17 44.935 ;
     RECT  1.19 47.545 121.17 50.375 ;
     RECT  1.19 52.985 121.17 55.815 ;
     RECT  1.19 58.425 121.17 61.255 ;
     RECT  1.19 63.865 121.17 66.695 ;
     RECT  1.19 69.305 121.17 72.135 ;
     RECT  1.19 74.745 121.17 77.575 ;
     RECT  1.19 80.185 121.17 83.015 ;
     RECT  1.19 85.625 121.17 88.455 ;
     RECT  1.19 91.065 121.17 93.895 ;
     RECT  1.19 96.505 121.17 99.335 ;
     RECT  1.19 101.945 121.17 104.775 ;
     RECT  1.19 107.385 121.17 110.215 ;
     RECT  1.19 112.825 121.17 115.655 ;
     RECT  1.19 118.265 121.17 121.095 ;
     RECT  1.19 123.705 121.17 126.535 ;
     RECT  1.19 129.145 121.17 131.975 ;
     RECT  1.19 134.585 121.17 137.415 ;
     RECT  1.19 140.025 121.17 142.855 ;
     RECT  1.19 145.465 121.17 148.295 ;
     RECT  1.19 150.905 121.17 153.735 ;
     RECT  1.19 156.345 121.17 159.175 ;
     RECT  1.19 161.785 121.17 164.615 ;
     RECT  1.19 167.225 121.17 170.055 ;
     RECT  1.19 172.665 121.17 175.495 ;
     RECT  1.19 178.105 121.17 180.935 ;
     RECT  1.19 183.545 121.17 186.375 ;
     RECT  1.19 188.985 121.17 191.815 ;
     RECT  1.19 194.425 121.17 197.255 ;
     RECT  1.19 199.865 121.17 202.695 ;
     RECT  1.19 205.305 121.17 208.135 ;
     RECT  1.19 210.745 121.17 213.575 ;
     RECT  1.19 216.185 121.17 219.015 ;
     RECT  1.19 221.625 121.17 224.455 ;
     RECT  1.19 227.065 121.17 229.895 ;
     RECT  1.19 232.505 121.17 235.335 ;
     RECT  1.19 237.945 121.17 239.55 ;
    LAYER pwell ;
     RECT  10.72 2.665 10.84 2.775 ;
     RECT  120.66 2.665 120.78 2.775 ;
     RECT  8.915 2.66 9.025 2.78 ;
     RECT  23.175 2.66 23.285 2.78 ;
     RECT  29.615 2.66 29.725 2.78 ;
     RECT  50.775 2.66 50.885 2.78 ;
     RECT  68.715 2.66 68.825 2.78 ;
     RECT  78.355 2.67 78.515 2.78 ;
     RECT  83.415 2.67 83.575 2.78 ;
     RECT  84.795 2.67 84.955 2.78 ;
     RECT  110.115 2.66 110.225 2.78 ;
     RECT  119.755 2.67 119.915 2.78 ;
     RECT  1.525 2.635 1.695 2.805 ;
     RECT  11.46 2.635 11.63 2.805 ;
     RECT  15.785 2.635 15.955 2.805 ;
     RECT  25.26 2.635 25.43 2.805 ;
     RECT  31.7 2.635 31.87 2.805 ;
     RECT  35.565 2.635 35.735 2.805 ;
     RECT  43.385 2.635 43.555 2.805 ;
     RECT  52.86 2.635 53.03 2.805 ;
     RECT  57.185 2.635 57.355 2.805 ;
     RECT  64.82 2.635 64.99 2.805 ;
     RECT  70.985 2.635 71.155 2.805 ;
     RECT  79.54 2.635 79.71 2.805 ;
     RECT  85.98 2.635 86.15 2.805 ;
     RECT  90.12 2.635 90.29 2.805 ;
     RECT  94.26 2.635 94.43 2.805 ;
     RECT  98.585 2.635 98.755 2.805 ;
     RECT  106.22 2.635 106.39 2.805 ;
     RECT  112.385 2.635 112.555 2.805 ;
     RECT  15.325 3.04 15.495 3.565 ;
     RECT  29.125 3.04 29.295 3.565 ;
     RECT  42.925 3.04 43.095 3.565 ;
     RECT  56.725 3.04 56.895 3.565 ;
     RECT  70.525 3.04 70.695 3.565 ;
     RECT  84.325 3.04 84.495 3.565 ;
     RECT  98.125 3.04 98.295 3.565 ;
     RECT  111.925 3.04 112.095 3.565 ;
     RECT  29.125 7.315 29.295 7.84 ;
     RECT  56.725 7.315 56.895 7.84 ;
     RECT  84.325 7.315 84.495 7.84 ;
     RECT  111.925 7.315 112.095 7.84 ;
     RECT  16.255 8.1 16.415 8.21 ;
     RECT  47.535 8.1 47.695 8.21 ;
     RECT  61.335 8.1 61.495 8.21 ;
     RECT  119.755 8.1 119.915 8.21 ;
     RECT  7.5 8.105 7.62 8.215 ;
     RECT  17.16 8.105 17.28 8.215 ;
     RECT  31.42 8.105 31.54 8.215 ;
     RECT  38.32 8.105 38.44 8.215 ;
     RECT  48.44 8.105 48.56 8.215 ;
     RECT  56.26 8.105 56.38 8.215 ;
     RECT  62.24 8.105 62.36 8.215 ;
     RECT  120.66 8.105 120.78 8.215 ;
     RECT  6.595 8.11 6.755 8.22 ;
     RECT  15.795 8.11 15.955 8.22 ;
     RECT  28.235 8.1 28.345 8.22 ;
     RECT  29.615 8.1 29.725 8.22 ;
     RECT  30.055 8.11 30.215 8.22 ;
     RECT  43.395 8.11 43.555 8.22 ;
     RECT  45.715 8.1 45.825 8.22 ;
     RECT  59.055 8.1 59.165 8.22 ;
     RECT  82.515 8.1 82.625 8.22 ;
     RECT  95.855 8.1 95.965 8.22 ;
     RECT  97.215 8.11 97.375 8.22 ;
     RECT  98.615 8.1 98.725 8.22 ;
     RECT  100.435 8.11 100.595 8.22 ;
     RECT  1.525 8.075 1.695 8.245 ;
     RECT  2.72 8.075 2.89 8.245 ;
     RECT  7.965 8.075 8.135 8.245 ;
     RECT  8.885 8.075 9.055 8.245 ;
     RECT  16.705 8.075 16.875 8.245 ;
     RECT  17.9 8.075 18.07 8.245 ;
     RECT  21.765 8.075 21.935 8.245 ;
     RECT  24.34 8.075 24.51 8.245 ;
     RECT  30.965 8.075 31.135 8.245 ;
     RECT  32.16 8.075 32.33 8.245 ;
     RECT  36.025 8.075 36.195 8.245 ;
     RECT  39.06 8.075 39.23 8.245 ;
     RECT  44.305 8.075 44.475 8.245 ;
     RECT  48.905 8.075 49.075 8.245 ;
     RECT  51.665 8.075 51.835 8.245 ;
     RECT  57.46 8.075 57.63 8.245 ;
     RECT  60.865 8.075 61.035 8.245 ;
     RECT  62.705 8.075 62.875 8.245 ;
     RECT  70.34 8.075 70.51 8.245 ;
     RECT  70.985 8.075 71.155 8.245 ;
     RECT  74.48 8.075 74.65 8.245 ;
     RECT  78.345 8.075 78.515 8.245 ;
     RECT  78.62 8.075 78.79 8.245 ;
     RECT  85.705 8.075 85.875 8.245 ;
     RECT  88.465 8.075 88.635 8.245 ;
     RECT  93.34 8.075 93.51 8.245 ;
     RECT  97.94 8.075 98.11 8.245 ;
     RECT  101.345 8.075 101.515 8.245 ;
     RECT  101.81 8.075 101.98 8.245 ;
     RECT  111.01 8.075 111.18 8.245 ;
     RECT  112.385 8.075 112.555 8.245 ;
     RECT  84.77 8.11 84.99 8.28 ;
     RECT  15.325 8.48 15.495 9.005 ;
     RECT  42.925 8.48 43.095 9.005 ;
     RECT  70.525 8.48 70.695 9.005 ;
     RECT  98.125 8.48 98.295 9.005 ;
     RECT  29.125 12.755 29.295 13.28 ;
     RECT  56.725 12.755 56.895 13.28 ;
     RECT  84.325 12.755 84.495 13.28 ;
     RECT  111.925 12.755 112.095 13.28 ;
     RECT  1.535 13.54 1.695 13.65 ;
     RECT  18.095 13.54 18.255 13.65 ;
     RECT  37.415 13.54 37.575 13.65 ;
     RECT  42.475 13.54 42.635 13.65 ;
     RECT  47.535 13.54 47.695 13.65 ;
     RECT  70.97 13.48 71.19 13.65 ;
     RECT  84.795 13.54 84.955 13.65 ;
     RECT  110.555 13.54 110.715 13.65 ;
     RECT  112.395 13.54 112.555 13.65 ;
     RECT  14.86 13.545 14.98 13.655 ;
     RECT  16.7 13.545 16.82 13.655 ;
     RECT  29.58 13.545 29.7 13.655 ;
     RECT  48.44 13.545 48.56 13.655 ;
     RECT  52.58 13.545 52.7 13.655 ;
     RECT  56.26 13.545 56.38 13.655 ;
     RECT  57.18 13.545 57.3 13.655 ;
     RECT  65.92 13.545 66.04 13.655 ;
     RECT  79.72 13.545 79.84 13.655 ;
     RECT  85.7 13.545 85.82 13.655 ;
     RECT  88 13.545 88.12 13.655 ;
     RECT  111.46 13.545 111.58 13.655 ;
     RECT  120.66 13.545 120.78 13.655 ;
     RECT  1.555 13.65 1.665 13.66 ;
     RECT  15.795 13.55 15.955 13.66 ;
     RECT  16.275 13.54 16.385 13.66 ;
     RECT  27.315 13.54 27.425 13.66 ;
     RECT  32.835 13.54 32.945 13.66 ;
     RECT  34.655 13.55 34.815 13.66 ;
     RECT  50.775 13.54 50.885 13.66 ;
     RECT  61.355 13.54 61.465 13.66 ;
     RECT  65.015 13.55 65.175 13.66 ;
     RECT  77.915 13.54 78.025 13.66 ;
     RECT  102.755 13.54 102.865 13.66 ;
     RECT  120.215 13.55 120.375 13.66 ;
     RECT  2.72 13.515 2.89 13.685 ;
     RECT  3.64 13.515 3.81 13.685 ;
     RECT  6.585 13.515 6.755 13.685 ;
     RECT  7.505 13.515 7.675 13.685 ;
     RECT  17.44 13.515 17.61 13.685 ;
     RECT  19.005 13.515 19.175 13.685 ;
     RECT  21.305 13.515 21.475 13.685 ;
     RECT  28.94 13.515 29.11 13.685 ;
     RECT  30.045 13.515 30.215 13.685 ;
     RECT  35.565 13.515 35.735 13.685 ;
     RECT  38.6 13.515 38.77 13.685 ;
     RECT  43.385 13.515 43.555 13.685 ;
     RECT  43.66 13.515 43.83 13.685 ;
     RECT  48.905 13.515 49.075 13.685 ;
     RECT  53.32 13.515 53.49 13.685 ;
     RECT  57.46 13.515 57.63 13.685 ;
     RECT  57.645 13.515 57.815 13.685 ;
     RECT  63.165 13.515 63.335 13.685 ;
     RECT  66.66 13.515 66.83 13.685 ;
     RECT  70.525 13.515 70.695 13.685 ;
     RECT  74.94 13.515 75.11 13.685 ;
     RECT  78.805 13.515 78.975 13.685 ;
     RECT  80.46 13.515 80.63 13.685 ;
     RECT  86.165 13.515 86.335 13.685 ;
     RECT  88.47 13.515 88.64 13.685 ;
     RECT  90.765 13.515 90.935 13.685 ;
     RECT  95.825 13.515 95.995 13.685 ;
     RECT  98.86 13.515 99.03 13.685 ;
     RECT  103.185 13.515 103.355 13.685 ;
     RECT  104.565 13.515 104.735 13.685 ;
     RECT  112.2 13.515 112.37 13.685 ;
     RECT  113.305 13.515 113.475 13.685 ;
     RECT  116.34 13.515 116.51 13.685 ;
     RECT  15.325 13.92 15.495 14.445 ;
     RECT  42.925 13.92 43.095 14.445 ;
     RECT  70.525 13.92 70.695 14.445 ;
     RECT  98.125 13.92 98.295 14.445 ;
     RECT  29.125 18.195 29.295 18.72 ;
     RECT  56.725 18.195 56.895 18.72 ;
     RECT  84.325 18.195 84.495 18.72 ;
     RECT  111.925 18.195 112.095 18.72 ;
     RECT  9.375 18.98 9.485 18.985 ;
     RECT  71.015 18.98 71.125 18.985 ;
     RECT  20.855 18.98 21.015 19.09 ;
     RECT  55.815 18.98 55.975 19.09 ;
     RECT  65.91 18.92 66.13 19.09 ;
     RECT  111.015 18.98 111.175 19.09 ;
     RECT  112.395 18.98 112.555 19.09 ;
     RECT  1.52 18.985 1.64 19.095 ;
     RECT  9.34 18.985 9.485 19.095 ;
     RECT  15.78 18.985 15.9 19.095 ;
     RECT  32.8 18.985 32.92 19.095 ;
     RECT  42.46 18.985 42.58 19.095 ;
     RECT  44.3 18.985 44.42 19.095 ;
     RECT  48.9 18.985 49.02 19.095 ;
     RECT  70.98 18.985 71.125 19.095 ;
     RECT  75.58 18.985 75.7 19.095 ;
     RECT  83.86 18.985 83.98 19.095 ;
     RECT  120.66 18.985 120.78 19.095 ;
     RECT  9.375 19.095 9.485 19.1 ;
     RECT  19.035 18.98 19.145 19.1 ;
     RECT  31.895 18.99 32.055 19.1 ;
     RECT  40.655 18.98 40.765 19.1 ;
     RECT  43.395 18.99 43.555 19.1 ;
     RECT  53.995 18.98 54.105 19.1 ;
     RECT  60.875 18.99 61.035 19.1 ;
     RECT  69.615 18.99 69.775 19.1 ;
     RECT  71.015 19.095 71.125 19.1 ;
     RECT  97.215 18.99 97.375 19.1 ;
     RECT  105.955 18.99 106.115 19.1 ;
     RECT  1.985 18.955 2.155 19.125 ;
     RECT  9.805 18.955 9.975 19.125 ;
     RECT  11.46 18.955 11.63 19.125 ;
     RECT  16.245 18.955 16.415 19.125 ;
     RECT  21.765 18.955 21.935 19.125 ;
     RECT  23.605 18.955 23.775 19.125 ;
     RECT  29.585 18.955 29.755 19.125 ;
     RECT  33.265 18.955 33.435 19.125 ;
     RECT  36.945 18.955 37.115 19.125 ;
     RECT  45.04 18.955 45.21 19.125 ;
     RECT  46.605 18.955 46.775 19.125 ;
     RECT  49.365 18.955 49.535 19.125 ;
     RECT  57 18.955 57.17 19.125 ;
     RECT  57.185 18.955 57.355 19.125 ;
     RECT  62.06 18.955 62.23 19.125 ;
     RECT  67.12 18.955 67.29 19.125 ;
     RECT  71.72 18.955 71.89 19.125 ;
     RECT  72.825 18.955 72.995 19.125 ;
     RECT  76.045 18.955 76.215 19.125 ;
     RECT  84.785 18.955 84.955 19.125 ;
     RECT  85.98 18.955 86.15 19.125 ;
     RECT  89.845 18.955 90.015 19.125 ;
     RECT  92.42 18.955 92.59 19.125 ;
     RECT  93.34 18.955 93.51 19.125 ;
     RECT  96.285 18.955 96.455 19.125 ;
     RECT  98.585 18.955 98.755 19.125 ;
     RECT  99.505 18.955 99.675 19.125 ;
     RECT  106.865 18.955 107.035 19.125 ;
     RECT  107.14 18.955 107.31 19.125 ;
     RECT  113.305 18.955 113.475 19.125 ;
     RECT  116.8 18.955 116.97 19.125 ;
     RECT  80.17 18.99 80.39 19.16 ;
     RECT  15.325 19.36 15.495 19.885 ;
     RECT  42.925 19.36 43.095 19.885 ;
     RECT  70.525 19.36 70.695 19.885 ;
     RECT  98.125 19.36 98.295 19.885 ;
     RECT  29.125 23.635 29.295 24.16 ;
     RECT  56.725 23.635 56.895 24.16 ;
     RECT  84.325 23.635 84.495 24.16 ;
     RECT  111.925 23.635 112.095 24.16 ;
     RECT  1.52 24.425 1.64 24.43 ;
     RECT  9.355 24.42 9.515 24.53 ;
     RECT  40.175 24.42 40.335 24.53 ;
     RECT  1.52 24.43 1.695 24.535 ;
     RECT  10.72 24.425 10.84 24.535 ;
     RECT  18.54 24.425 18.66 24.535 ;
     RECT  29.58 24.425 29.7 24.535 ;
     RECT  35.1 24.425 35.22 24.535 ;
     RECT  52.58 24.425 52.7 24.535 ;
     RECT  56.26 24.425 56.38 24.535 ;
     RECT  59.94 24.425 60.06 24.535 ;
     RECT  66.38 24.425 66.5 24.535 ;
     RECT  73.74 24.425 73.86 24.535 ;
     RECT  83.86 24.425 83.98 24.535 ;
     RECT  93.52 24.425 93.64 24.535 ;
     RECT  98.12 24.425 98.24 24.535 ;
     RECT  120.66 24.425 120.78 24.535 ;
     RECT  1.535 24.535 1.695 24.54 ;
     RECT  9.815 24.43 9.975 24.54 ;
     RECT  15.815 24.42 15.925 24.54 ;
     RECT  17.635 24.43 17.795 24.54 ;
     RECT  33.295 24.42 33.405 24.54 ;
     RECT  51.675 24.43 51.835 24.54 ;
     RECT  54.455 24.42 54.565 24.54 ;
     RECT  57.215 24.42 57.325 24.54 ;
     RECT  59.035 24.42 59.195 24.54 ;
     RECT  64.575 24.42 64.685 24.54 ;
     RECT  68.715 24.42 68.825 24.54 ;
     RECT  71.015 24.42 71.125 24.54 ;
     RECT  72.835 24.43 72.995 24.54 ;
     RECT  88.955 24.42 89.065 24.54 ;
     RECT  98.615 24.42 98.725 24.54 ;
     RECT  100.435 24.43 100.595 24.54 ;
     RECT  1.985 24.395 2.155 24.565 ;
     RECT  2.445 24.395 2.615 24.565 ;
     RECT  10.54 24.395 10.71 24.565 ;
     RECT  11.46 24.395 11.63 24.565 ;
     RECT  14.405 24.395 14.575 24.565 ;
     RECT  19.28 24.395 19.45 24.565 ;
     RECT  21.765 24.395 21.935 24.565 ;
     RECT  23.15 24.395 23.32 24.565 ;
     RECT  30.32 24.395 30.49 24.565 ;
     RECT  34.19 24.395 34.36 24.565 ;
     RECT  35.565 24.395 35.735 24.565 ;
     RECT  41.085 24.395 41.255 24.565 ;
     RECT  43.385 24.395 43.555 24.565 ;
     RECT  50.56 24.395 50.73 24.565 ;
     RECT  53.32 24.395 53.49 24.565 ;
     RECT  60.405 24.395 60.575 24.565 ;
     RECT  60.68 24.395 60.85 24.565 ;
     RECT  66.845 24.395 67.015 24.565 ;
     RECT  74.205 24.395 74.375 24.565 ;
     RECT  74.48 24.395 74.65 24.565 ;
     RECT  78.345 24.395 78.515 24.565 ;
     RECT  85.06 24.395 85.23 24.565 ;
     RECT  85.71 24.395 85.88 24.565 ;
     RECT  90.765 24.395 90.935 24.565 ;
     RECT  94.26 24.395 94.43 24.565 ;
     RECT  98.86 24.395 99.03 24.565 ;
     RECT  101.345 24.395 101.515 24.565 ;
     RECT  102.725 24.395 102.895 24.565 ;
     RECT  111.01 24.395 111.18 24.565 ;
     RECT  112.66 24.395 112.83 24.565 ;
     RECT  116.8 24.395 116.97 24.565 ;
     RECT  15.325 24.8 15.495 25.325 ;
     RECT  42.925 24.8 43.095 25.325 ;
     RECT  70.525 24.8 70.695 25.325 ;
     RECT  98.125 24.8 98.295 25.325 ;
     RECT  29.125 29.075 29.295 29.6 ;
     RECT  56.725 29.075 56.895 29.6 ;
     RECT  84.325 29.075 84.495 29.6 ;
     RECT  111.925 29.075 112.095 29.6 ;
     RECT  1.555 29.86 1.665 29.865 ;
     RECT  55.355 29.86 55.515 29.97 ;
     RECT  64.99 29.8 65.21 29.97 ;
     RECT  70.97 29.8 71.19 29.97 ;
     RECT  92.155 29.86 92.315 29.97 ;
     RECT  112.395 29.86 112.555 29.97 ;
     RECT  1.52 29.865 1.665 29.975 ;
     RECT  3.36 29.865 3.48 29.975 ;
     RECT  33.72 29.865 33.84 29.975 ;
     RECT  38.32 29.865 38.44 29.975 ;
     RECT  45.22 29.865 45.34 29.975 ;
     RECT  49.82 29.865 49.94 29.975 ;
     RECT  56.26 29.865 56.38 29.975 ;
     RECT  59.02 29.865 59.14 29.975 ;
     RECT  75.58 29.865 75.7 29.975 ;
     RECT  99.5 29.865 99.62 29.975 ;
     RECT  120.66 29.865 120.78 29.975 ;
     RECT  1.555 29.975 1.665 29.98 ;
     RECT  23.175 29.86 23.285 29.98 ;
     RECT  28.215 29.87 28.375 29.98 ;
     RECT  43.415 29.86 43.525 29.98 ;
     RECT  57.215 29.86 57.325 29.98 ;
     RECT  68.715 29.86 68.825 29.98 ;
     RECT  74.675 29.87 74.835 29.98 ;
     RECT  90.335 29.86 90.445 29.98 ;
     RECT  98.595 29.87 98.755 29.98 ;
     RECT  2.26 29.835 2.43 30.005 ;
     RECT  4.1 29.835 4.27 30.005 ;
     RECT  6.125 29.835 6.295 30.005 ;
     RECT  7.965 29.835 8.135 30.005 ;
     RECT  15.785 29.835 15.955 30.005 ;
     RECT  24.34 29.835 24.51 30.005 ;
     RECT  25.26 29.835 25.43 30.005 ;
     RECT  29.125 29.835 29.295 30.005 ;
     RECT  29.86 29.835 30.03 30.005 ;
     RECT  34.19 29.835 34.36 30.005 ;
     RECT  39.06 29.835 39.23 30.005 ;
     RECT  44.305 29.835 44.475 30.005 ;
     RECT  45.96 29.835 46.13 30.005 ;
     RECT  50.285 29.835 50.455 30.005 ;
     RECT  57.645 29.835 57.815 30.005 ;
     RECT  59.485 29.835 59.655 30.005 ;
     RECT  67.12 29.835 67.29 30.005 ;
     RECT  71.905 29.835 72.075 30.005 ;
     RECT  76.045 29.835 76.215 30.005 ;
     RECT  79.54 29.835 79.71 30.005 ;
     RECT  83.405 29.835 83.575 30.005 ;
     RECT  84.785 29.835 84.955 30.005 ;
     RECT  88.01 29.835 88.18 30.005 ;
     RECT  90.765 29.835 90.935 30.005 ;
     RECT  93.34 29.835 93.51 30.005 ;
     RECT  97.205 29.835 97.375 30.005 ;
     RECT  100.24 29.835 100.41 30.005 ;
     RECT  104.105 29.835 104.275 30.005 ;
     RECT  104.565 29.835 104.735 30.005 ;
     RECT  108.06 29.835 108.23 30.005 ;
     RECT  111.465 29.835 111.635 30.005 ;
     RECT  113.305 29.835 113.475 30.005 ;
     RECT  51.65 29.87 51.87 30.04 ;
     RECT  15.325 30.24 15.495 30.765 ;
     RECT  42.925 30.24 43.095 30.765 ;
     RECT  70.525 30.24 70.695 30.765 ;
     RECT  98.125 30.24 98.295 30.765 ;
     RECT  29.125 34.515 29.295 35.04 ;
     RECT  56.725 34.515 56.895 35.04 ;
     RECT  84.325 34.515 84.495 35.04 ;
     RECT  111.925 34.515 112.095 35.04 ;
     RECT  28.215 35.3 28.375 35.41 ;
     RECT  36.955 35.3 37.115 35.41 ;
     RECT  43.37 35.24 43.59 35.41 ;
     RECT  65.015 35.3 65.175 35.41 ;
     RECT  112.395 35.3 112.555 35.41 ;
     RECT  3.36 35.305 3.48 35.415 ;
     RECT  14.86 35.305 14.98 35.415 ;
     RECT  20.38 35.305 20.5 35.415 ;
     RECT  37.86 35.305 37.98 35.415 ;
     RECT  42.46 35.305 42.58 35.415 ;
     RECT  53.04 35.305 53.16 35.415 ;
     RECT  65.92 35.305 66.04 35.415 ;
     RECT  70.06 35.305 70.18 35.415 ;
     RECT  83.86 35.305 83.98 35.415 ;
     RECT  98.58 35.305 98.7 35.415 ;
     RECT  107.32 35.305 107.44 35.415 ;
     RECT  120.66 35.305 120.78 35.415 ;
     RECT  7.995 35.3 8.105 35.42 ;
     RECT  9.815 35.31 9.975 35.42 ;
     RECT  19.955 35.3 20.065 35.42 ;
     RECT  35.595 35.3 35.705 35.42 ;
     RECT  37.415 35.31 37.575 35.42 ;
     RECT  51.235 35.3 51.345 35.42 ;
     RECT  71.015 35.3 71.125 35.42 ;
     RECT  72.835 35.31 72.995 35.42 ;
     RECT  82.055 35.3 82.165 35.42 ;
     RECT  97.215 35.31 97.375 35.42 ;
     RECT  106.415 35.31 106.575 35.42 ;
     RECT  119.315 35.3 119.425 35.42 ;
     RECT  1.525 35.275 1.695 35.445 ;
     RECT  4.1 35.275 4.27 35.445 ;
     RECT  9.16 35.275 9.33 35.445 ;
     RECT  11 35.275 11.17 35.445 ;
     RECT  13.025 35.275 13.195 35.445 ;
     RECT  16.06 35.275 16.23 35.445 ;
     RECT  20.845 35.275 21.015 35.445 ;
     RECT  22.04 35.275 22.21 35.445 ;
     RECT  25.905 35.275 26.075 35.445 ;
     RECT  29.585 35.275 29.755 35.445 ;
     RECT  38.325 35.275 38.495 35.445 ;
     RECT  38.6 35.275 38.77 35.445 ;
     RECT  47.34 35.275 47.51 35.445 ;
     RECT  49.365 35.275 49.535 35.445 ;
     RECT  53.505 35.275 53.675 35.445 ;
     RECT  57.46 35.275 57.63 35.445 ;
     RECT  62.705 35.275 62.875 35.445 ;
     RECT  66.385 35.275 66.555 35.445 ;
     RECT  73.745 35.275 73.915 35.445 ;
     RECT  74.02 35.275 74.19 35.445 ;
     RECT  78.16 35.275 78.33 35.445 ;
     RECT  83.68 35.275 83.85 35.445 ;
     RECT  84.785 35.275 84.955 35.445 ;
     RECT  87.545 35.275 87.715 35.445 ;
     RECT  92.145 35.275 92.315 35.445 ;
     RECT  99.045 35.275 99.215 35.445 ;
     RECT  99.78 35.275 99.95 35.445 ;
     RECT  103.92 35.275 104.09 35.445 ;
     RECT  107.785 35.275 107.955 35.445 ;
     RECT  108.06 35.275 108.23 35.445 ;
     RECT  113.305 35.275 113.475 35.445 ;
     RECT  115.42 35.275 115.59 35.445 ;
     RECT  45.67 35.31 45.89 35.48 ;
     RECT  61.31 35.31 61.53 35.48 ;
     RECT  15.325 35.68 15.495 36.205 ;
     RECT  42.925 35.68 43.095 36.205 ;
     RECT  70.525 35.68 70.695 36.205 ;
     RECT  98.125 35.68 98.295 36.205 ;
     RECT  29.125 39.955 29.295 40.48 ;
     RECT  56.725 39.955 56.895 40.48 ;
     RECT  84.325 39.955 84.495 40.48 ;
     RECT  111.925 39.955 112.095 40.48 ;
     RECT  70.075 40.74 70.235 40.745 ;
     RECT  111.465 40.715 111.635 40.745 ;
     RECT  1.52 40.745 1.64 40.75 ;
     RECT  70.06 40.745 70.235 40.85 ;
     RECT  93.075 40.74 93.235 40.85 ;
     RECT  110.555 40.74 110.715 40.85 ;
     RECT  120.215 40.74 120.375 40.85 ;
     RECT  1.52 40.75 1.695 40.855 ;
     RECT  2.44 40.745 2.56 40.855 ;
     RECT  34.18 40.745 34.3 40.855 ;
     RECT  58.1 40.745 58.22 40.855 ;
     RECT  64.54 40.745 64.66 40.855 ;
     RECT  70.06 40.85 70.18 40.855 ;
     RECT  111 40.745 111.12 40.855 ;
     RECT  111.46 40.745 111.635 40.855 ;
     RECT  115.6 40.745 115.72 40.855 ;
     RECT  1.535 40.855 1.695 40.86 ;
     RECT  7.055 40.75 7.215 40.86 ;
     RECT  68.255 40.74 68.365 40.86 ;
     RECT  69.155 40.75 69.315 40.86 ;
     RECT  82.515 40.74 82.625 40.86 ;
     RECT  98.595 40.75 98.755 40.86 ;
     RECT  109.195 40.74 109.305 40.86 ;
     RECT  1.985 40.715 2.155 40.885 ;
     RECT  3.18 40.715 3.35 40.885 ;
     RECT  7.965 40.715 8.135 40.885 ;
     RECT  9.345 40.715 9.515 40.885 ;
     RECT  16.06 40.715 16.23 40.885 ;
     RECT  16.98 40.715 17.15 40.885 ;
     RECT  20.2 40.715 20.37 40.885 ;
     RECT  21.12 40.715 21.29 40.885 ;
     RECT  24.065 40.715 24.235 40.885 ;
     RECT  25.26 40.715 25.43 40.885 ;
     RECT  29.59 40.715 29.76 40.885 ;
     RECT  31.425 40.715 31.595 40.885 ;
     RECT  34.645 40.715 34.815 40.885 ;
     RECT  39.06 40.715 39.23 40.885 ;
     RECT  42.005 40.715 42.175 40.885 ;
     RECT  43.385 40.715 43.555 40.885 ;
     RECT  49.365 40.715 49.535 40.885 ;
     RECT  53.32 40.715 53.49 40.885 ;
     RECT  57.185 40.715 57.355 40.885 ;
     RECT  58.565 40.715 58.735 40.885 ;
     RECT  65.28 40.715 65.45 40.885 ;
     RECT  70.985 40.715 71.155 40.885 ;
     RECT  78.62 40.715 78.79 40.885 ;
     RECT  80.185 40.715 80.355 40.885 ;
     RECT  85.06 40.715 85.23 40.885 ;
     RECT  87.545 40.715 87.715 40.885 ;
     RECT  89.2 40.715 89.37 40.885 ;
     RECT  90.765 40.715 90.935 40.885 ;
     RECT  93.985 40.715 94.155 40.885 ;
     RECT  99.505 40.715 99.675 40.885 ;
     RECT  103.185 40.715 103.355 40.885 ;
     RECT  111.465 40.855 111.635 40.885 ;
     RECT  112.385 40.715 112.555 40.885 ;
     RECT  116.34 40.715 116.51 40.885 ;
     RECT  15.325 41.12 15.495 41.645 ;
     RECT  42.925 41.12 43.095 41.645 ;
     RECT  70.525 41.12 70.695 41.645 ;
     RECT  98.125 41.12 98.295 41.645 ;
     RECT  29.125 45.395 29.295 45.92 ;
     RECT  56.725 45.395 56.895 45.92 ;
     RECT  84.325 45.395 84.495 45.92 ;
     RECT  111.925 45.395 112.095 45.92 ;
     RECT  1.535 46.18 1.695 46.185 ;
     RECT  16.715 46.18 16.875 46.185 ;
     RECT  65.925 46.155 66.095 46.185 ;
     RECT  1.52 46.185 1.695 46.29 ;
     RECT  16.7 46.185 16.875 46.29 ;
     RECT  60.39 46.12 60.61 46.29 ;
     RECT  73.295 46.18 73.455 46.29 ;
     RECT  119.755 46.18 119.915 46.29 ;
     RECT  1.52 46.29 1.64 46.295 ;
     RECT  2.44 46.185 2.56 46.295 ;
     RECT  16.7 46.29 16.82 46.295 ;
     RECT  35.1 46.185 35.22 46.295 ;
     RECT  52.58 46.185 52.7 46.295 ;
     RECT  56.26 46.185 56.38 46.295 ;
     RECT  60.86 46.185 60.98 46.295 ;
     RECT  65.46 46.185 65.58 46.295 ;
     RECT  65.92 46.185 66.095 46.295 ;
     RECT  74.2 46.185 74.32 46.295 ;
     RECT  85.24 46.185 85.36 46.295 ;
     RECT  120.66 46.185 120.78 46.295 ;
     RECT  9.375 46.18 9.485 46.3 ;
     RECT  15.795 46.19 15.955 46.3 ;
     RECT  34.195 46.19 34.355 46.3 ;
     RECT  43.415 46.18 43.525 46.3 ;
     RECT  54.455 46.18 54.565 46.3 ;
     RECT  64.115 46.18 64.225 46.3 ;
     RECT  78.355 46.19 78.515 46.3 ;
     RECT  83.435 46.18 83.545 46.3 ;
     RECT  97.215 46.19 97.375 46.3 ;
     RECT  98.615 46.18 98.725 46.3 ;
     RECT  100.435 46.19 100.595 46.3 ;
     RECT  112.855 46.19 113.015 46.3 ;
     RECT  1.985 46.155 2.155 46.325 ;
     RECT  3.18 46.155 3.35 46.325 ;
     RECT  7.045 46.155 7.215 46.325 ;
     RECT  11.46 46.155 11.63 46.325 ;
     RECT  17.165 46.155 17.335 46.325 ;
     RECT  17.9 46.155 18.07 46.325 ;
     RECT  21.765 46.155 21.935 46.325 ;
     RECT  24.525 46.155 24.695 46.325 ;
     RECT  29.585 46.155 29.755 46.325 ;
     RECT  35.565 46.155 35.735 46.325 ;
     RECT  36.95 46.155 37.12 46.325 ;
     RECT  42.925 46.155 43.095 46.325 ;
     RECT  45.225 46.155 45.395 46.325 ;
     RECT  50.56 46.155 50.73 46.325 ;
     RECT  53.045 46.155 53.215 46.325 ;
     RECT  61.6 46.155 61.77 46.325 ;
     RECT  65.925 46.295 66.095 46.325 ;
     RECT  66.66 46.155 66.83 46.325 ;
     RECT  70.985 46.155 71.155 46.325 ;
     RECT  74.665 46.155 74.835 46.325 ;
     RECT  79.54 46.155 79.71 46.325 ;
     RECT  82.03 46.155 82.2 46.325 ;
     RECT  85.06 46.155 85.23 46.325 ;
     RECT  85.705 46.155 85.875 46.325 ;
     RECT  88.925 46.155 89.095 46.325 ;
     RECT  93.34 46.155 93.51 46.325 ;
     RECT  96.56 46.155 96.73 46.325 ;
     RECT  100.7 46.155 100.87 46.325 ;
     RECT  101.62 46.155 101.79 46.325 ;
     RECT  104.84 46.155 105.01 46.325 ;
     RECT  105.485 46.155 105.655 46.325 ;
     RECT  108.705 46.155 108.875 46.325 ;
     RECT  112.385 46.155 112.555 46.325 ;
     RECT  113.765 46.155 113.935 46.325 ;
     RECT  57.17 46.19 57.39 46.36 ;
     RECT  15.325 46.56 15.495 47.085 ;
     RECT  42.925 46.56 43.095 47.085 ;
     RECT  70.525 46.56 70.695 47.085 ;
     RECT  98.125 46.56 98.295 47.085 ;
     RECT  29.125 50.835 29.295 51.36 ;
     RECT  56.725 50.835 56.895 51.36 ;
     RECT  84.325 50.835 84.495 51.36 ;
     RECT  111.925 50.835 112.095 51.36 ;
     RECT  1.535 51.62 1.695 51.73 ;
     RECT  28.215 51.62 28.375 51.73 ;
     RECT  29.11 51.56 29.33 51.73 ;
     RECT  41.555 51.62 41.715 51.73 ;
     RECT  72.375 51.62 72.535 51.73 ;
     RECT  82.955 51.62 83.115 51.73 ;
     RECT  112.395 51.62 112.555 51.73 ;
     RECT  3.36 51.625 3.48 51.735 ;
     RECT  36.94 51.625 37.06 51.735 ;
     RECT  46.6 51.625 46.72 51.735 ;
     RECT  83.86 51.625 83.98 51.735 ;
     RECT  99.5 51.625 99.62 51.735 ;
     RECT  111.46 51.625 111.58 51.735 ;
     RECT  113.3 51.625 113.42 51.735 ;
     RECT  120.66 51.625 120.78 51.735 ;
     RECT  1.555 51.73 1.665 51.74 ;
     RECT  15.795 51.63 15.955 51.74 ;
     RECT  26.395 51.62 26.505 51.74 ;
     RECT  32.815 51.63 32.975 51.74 ;
     RECT  35.135 51.62 35.245 51.74 ;
     RECT  53.055 51.63 53.215 51.74 ;
     RECT  54.915 51.62 55.025 51.74 ;
     RECT  61.355 51.62 61.465 51.74 ;
     RECT  70.995 51.63 71.155 51.74 ;
     RECT  96.315 51.62 96.425 51.74 ;
     RECT  98.595 51.63 98.755 51.74 ;
     RECT  103.675 51.62 103.785 51.74 ;
     RECT  107.335 51.63 107.495 51.74 ;
     RECT  109.655 51.62 109.765 51.74 ;
     RECT  119.755 51.63 119.915 51.74 ;
     RECT  2.445 51.595 2.615 51.765 ;
     RECT  4.1 51.595 4.27 51.765 ;
     RECT  7.965 51.595 8.135 51.765 ;
     RECT  9.805 51.595 9.975 51.765 ;
     RECT  16.98 51.595 17.15 51.765 ;
     RECT  19.005 51.595 19.175 51.765 ;
     RECT  21.12 51.595 21.29 51.765 ;
     RECT  25.26 51.595 25.43 51.765 ;
     RECT  29.86 51.595 30.03 51.765 ;
     RECT  33.72 51.595 33.9 51.765 ;
     RECT  35.565 51.595 35.735 51.765 ;
     RECT  37.68 51.595 37.85 51.765 ;
     RECT  42.74 51.595 42.91 51.765 ;
     RECT  43.385 51.595 43.555 51.765 ;
     RECT  47.34 51.595 47.51 51.765 ;
     RECT  53.965 51.595 54.135 51.765 ;
     RECT  57.46 51.595 57.63 51.765 ;
     RECT  63.165 51.595 63.335 51.765 ;
     RECT  64.36 51.595 64.53 51.765 ;
     RECT  68.5 51.595 68.67 51.765 ;
     RECT  71.905 51.595 72.075 51.765 ;
     RECT  73.285 51.595 73.455 51.765 ;
     RECT  79.265 51.595 79.435 51.765 ;
     RECT  84.785 51.595 84.955 51.765 ;
     RECT  86.625 51.595 86.795 51.765 ;
     RECT  92.145 51.595 92.315 51.765 ;
     RECT  99.78 51.595 99.95 51.765 ;
     RECT  99.965 51.595 100.135 51.765 ;
     RECT  105.76 51.595 105.93 51.765 ;
     RECT  108.245 51.595 108.415 51.765 ;
     RECT  113.765 51.595 113.935 51.765 ;
     RECT  115.88 51.595 116.05 51.765 ;
     RECT  51.19 51.63 51.41 51.8 ;
     RECT  15.325 52 15.495 52.525 ;
     RECT  42.925 52 43.095 52.525 ;
     RECT  70.525 52 70.695 52.525 ;
     RECT  98.125 52 98.295 52.525 ;
     RECT  29.125 56.275 29.295 56.8 ;
     RECT  56.725 56.275 56.895 56.8 ;
     RECT  84.325 56.275 84.495 56.8 ;
     RECT  111.925 56.275 112.095 56.8 ;
     RECT  1.555 57.06 1.665 57.07 ;
     RECT  7.515 57.06 7.675 57.17 ;
     RECT  57.195 57.06 57.355 57.17 ;
     RECT  63.61 57 63.83 57.17 ;
     RECT  64.095 57.06 64.255 57.17 ;
     RECT  79.275 57.06 79.435 57.17 ;
     RECT  84.795 57.06 84.955 57.17 ;
     RECT  2.44 57.065 2.56 57.175 ;
     RECT  8.42 57.065 8.54 57.175 ;
     RECT  15.78 57.065 15.9 57.175 ;
     RECT  17.16 57.065 17.28 57.175 ;
     RECT  29.58 57.065 29.7 57.175 ;
     RECT  44.3 57.065 44.42 57.175 ;
     RECT  56.26 57.065 56.38 57.175 ;
     RECT  65 57.065 65.12 57.175 ;
     RECT  76.04 57.065 76.16 57.175 ;
     RECT  88 57.065 88.12 57.175 ;
     RECT  89.84 57.065 89.96 57.175 ;
     RECT  100.42 57.065 100.54 57.175 ;
     RECT  101.8 57.065 101.92 57.175 ;
     RECT  112.38 57.065 112.5 57.175 ;
     RECT  1.535 57.07 1.695 57.18 ;
     RECT  14.415 57.07 14.575 57.18 ;
     RECT  34.655 57.07 34.815 57.18 ;
     RECT  43.395 57.07 43.555 57.18 ;
     RECT  62.275 57.06 62.385 57.18 ;
     RECT  70.995 57.07 71.155 57.18 ;
     RECT  98.615 57.06 98.725 57.18 ;
     RECT  2.905 57.035 3.075 57.205 ;
     RECT  3.64 57.035 3.81 57.205 ;
     RECT  8.885 57.035 9.055 57.205 ;
     RECT  10.54 57.035 10.71 57.205 ;
     RECT  16.245 57.035 16.415 57.205 ;
     RECT  17.9 57.035 18.07 57.205 ;
     RECT  21.765 57.035 21.935 57.205 ;
     RECT  23.605 57.035 23.775 57.205 ;
     RECT  30.32 57.035 30.49 57.205 ;
     RECT  33.26 57.035 33.43 57.205 ;
     RECT  34.19 57.035 34.36 57.205 ;
     RECT  35.565 57.035 35.735 57.205 ;
     RECT  44.58 57.035 44.75 57.205 ;
     RECT  44.765 57.035 44.935 57.205 ;
     RECT  48.72 57.035 48.89 57.205 ;
     RECT  52.125 57.035 52.295 57.205 ;
     RECT  58.38 57.035 58.55 57.205 ;
     RECT  59.76 57.035 59.93 57.205 ;
     RECT  65.465 57.035 65.635 57.205 ;
     RECT  67.305 57.035 67.475 57.205 ;
     RECT  72.18 57.035 72.35 57.205 ;
     RECT  75.4 57.035 75.57 57.205 ;
     RECT  76.78 57.035 76.95 57.205 ;
     RECT  80.46 57.035 80.63 57.205 ;
     RECT  80.645 57.035 80.815 57.205 ;
     RECT  85.98 57.035 86.15 57.205 ;
     RECT  88.47 57.035 88.64 57.205 ;
     RECT  90.305 57.035 90.475 57.205 ;
     RECT  90.765 57.035 90.935 57.205 ;
     RECT  93.525 57.035 93.695 57.205 ;
     RECT  100.885 57.035 101.055 57.205 ;
     RECT  102.265 57.035 102.435 57.205 ;
     RECT  108.245 57.035 108.415 57.205 ;
     RECT  111.465 57.035 111.635 57.205 ;
     RECT  113.12 57.035 113.29 57.205 ;
     RECT  117.26 57.035 117.43 57.205 ;
     RECT  52.57 57.07 52.79 57.24 ;
     RECT  15.325 57.44 15.495 57.965 ;
     RECT  42.925 57.44 43.095 57.965 ;
     RECT  70.525 57.44 70.695 57.965 ;
     RECT  98.125 57.44 98.295 57.965 ;
     RECT  29.125 61.715 29.295 62.24 ;
     RECT  56.725 61.715 56.895 62.24 ;
     RECT  84.325 61.715 84.495 62.24 ;
     RECT  111.925 61.715 112.095 62.24 ;
     RECT  1.555 62.5 1.665 62.505 ;
     RECT  23.615 62.5 23.775 62.61 ;
     RECT  55.815 62.5 55.975 62.61 ;
     RECT  65.475 62.5 65.635 62.61 ;
     RECT  76.055 62.5 76.215 62.61 ;
     RECT  93.075 62.5 93.235 62.61 ;
     RECT  119.755 62.5 119.915 62.61 ;
     RECT  1.52 62.505 1.665 62.615 ;
     RECT  3.36 62.505 3.48 62.615 ;
     RECT  7.96 62.505 8.08 62.615 ;
     RECT  10.26 62.505 10.38 62.615 ;
     RECT  14.86 62.505 14.98 62.615 ;
     RECT  15.78 62.505 15.9 62.615 ;
     RECT  24.52 62.505 24.64 62.615 ;
     RECT  38.78 62.505 38.9 62.615 ;
     RECT  66.38 62.505 66.5 62.615 ;
     RECT  84.32 62.505 84.44 62.615 ;
     RECT  93.98 62.505 94.1 62.615 ;
     RECT  120.66 62.505 120.78 62.615 ;
     RECT  1.555 62.615 1.665 62.62 ;
     RECT  9.355 62.51 9.515 62.62 ;
     RECT  60.435 62.5 60.545 62.62 ;
     RECT  62.255 62.51 62.415 62.62 ;
     RECT  71.015 62.5 71.125 62.62 ;
     RECT  72.835 62.51 72.995 62.62 ;
     RECT  74.235 62.5 74.345 62.62 ;
     RECT  83.415 62.51 83.575 62.62 ;
     RECT  96.315 62.5 96.425 62.62 ;
     RECT  98.615 62.5 98.725 62.62 ;
     RECT  102.755 62.5 102.865 62.62 ;
     RECT  1.985 62.475 2.155 62.645 ;
     RECT  4.1 62.475 4.27 62.645 ;
     RECT  8.425 62.475 8.595 62.645 ;
     RECT  11 62.475 11.17 62.645 ;
     RECT  16.06 62.475 16.23 62.645 ;
     RECT  16.245 62.475 16.415 62.645 ;
     RECT  20.2 62.475 20.37 62.645 ;
     RECT  24.34 62.475 24.51 62.645 ;
     RECT  25.26 62.475 25.43 62.645 ;
     RECT  28.205 62.475 28.375 62.645 ;
     RECT  29.59 62.475 29.76 62.645 ;
     RECT  31.425 62.475 31.595 62.645 ;
     RECT  35.565 62.475 35.735 62.645 ;
     RECT  39.245 62.475 39.415 62.645 ;
     RECT  43.385 62.475 43.555 62.645 ;
     RECT  48.445 62.475 48.615 62.645 ;
     RECT  53.045 62.475 53.215 62.645 ;
     RECT  57.46 62.475 57.63 62.645 ;
     RECT  61.6 62.475 61.77 62.645 ;
     RECT  63.165 62.475 63.335 62.645 ;
     RECT  66.845 62.475 67.015 62.645 ;
     RECT  73.745 62.475 73.915 62.645 ;
     RECT  76.965 62.475 77.135 62.645 ;
     RECT  84.785 62.475 84.955 62.645 ;
     RECT  85.06 62.475 85.23 62.645 ;
     RECT  89.2 62.475 89.37 62.645 ;
     RECT  92.42 62.475 92.59 62.645 ;
     RECT  94.72 62.475 94.89 62.645 ;
     RECT  98.86 62.475 99.03 62.645 ;
     RECT  100.425 62.475 100.595 62.645 ;
     RECT  104.565 62.475 104.735 62.645 ;
     RECT  107.785 62.475 107.955 62.645 ;
     RECT  112.385 62.475 112.555 62.645 ;
     RECT  117.26 62.475 117.43 62.645 ;
     RECT  15.325 62.88 15.495 63.405 ;
     RECT  42.925 62.88 43.095 63.405 ;
     RECT  70.525 62.88 70.695 63.405 ;
     RECT  98.125 62.88 98.295 63.405 ;
     RECT  29.125 67.155 29.295 67.68 ;
     RECT  56.725 67.155 56.895 67.68 ;
     RECT  84.325 67.155 84.495 67.68 ;
     RECT  111.925 67.155 112.095 67.68 ;
     RECT  59.025 67.915 59.195 67.945 ;
     RECT  1.555 67.94 1.665 67.95 ;
     RECT  18.555 67.94 18.715 68.05 ;
     RECT  46.155 67.94 46.315 68.05 ;
     RECT  84.795 67.94 84.955 68.05 ;
     RECT  110.555 67.94 110.715 68.05 ;
     RECT  2.44 67.945 2.56 68.055 ;
     RECT  3.36 67.945 3.48 68.055 ;
     RECT  28.66 67.945 28.78 68.055 ;
     RECT  29.58 67.945 29.7 68.055 ;
     RECT  47.06 67.945 47.18 68.055 ;
     RECT  54.42 67.945 54.54 68.055 ;
     RECT  59.02 67.945 59.195 68.055 ;
     RECT  83.86 67.945 83.98 68.055 ;
     RECT  111.46 67.945 111.58 68.055 ;
     RECT  116.52 67.945 116.64 68.055 ;
     RECT  120.66 67.945 120.78 68.055 ;
     RECT  1.535 67.95 1.695 68.06 ;
     RECT  26.855 67.94 26.965 68.06 ;
     RECT  44.335 67.94 44.445 68.06 ;
     RECT  52.615 67.94 52.725 68.06 ;
     RECT  54.915 67.94 55.025 68.06 ;
     RECT  57.215 67.94 57.325 68.06 ;
     RECT  97.215 67.95 97.375 68.06 ;
     RECT  3.18 67.915 3.35 68.085 ;
     RECT  3.825 67.915 3.995 68.085 ;
     RECT  7.045 67.915 7.215 68.085 ;
     RECT  11.185 67.915 11.355 68.085 ;
     RECT  16.06 67.915 16.23 68.085 ;
     RECT  19.465 67.915 19.635 68.085 ;
     RECT  20.2 67.915 20.37 68.085 ;
     RECT  24.34 67.915 24.51 68.085 ;
     RECT  28.205 67.915 28.375 68.085 ;
     RECT  30.32 67.915 30.49 68.085 ;
     RECT  34.19 67.915 34.36 68.085 ;
     RECT  35.565 67.915 35.735 68.085 ;
     RECT  43.385 67.915 43.555 68.085 ;
     RECT  47.525 67.915 47.695 68.085 ;
     RECT  55.16 67.915 55.33 68.085 ;
     RECT  59.025 68.055 59.195 68.085 ;
     RECT  59.485 67.915 59.655 68.085 ;
     RECT  66.66 67.915 66.83 68.085 ;
     RECT  69.145 67.915 69.315 68.085 ;
     RECT  70.985 67.915 71.155 68.085 ;
     RECT  76.78 67.915 76.95 68.085 ;
     RECT  78.345 67.915 78.515 68.085 ;
     RECT  80.645 67.915 80.815 68.085 ;
     RECT  85.705 67.915 85.875 68.085 ;
     RECT  93.34 67.915 93.51 68.085 ;
     RECT  94.905 67.915 95.075 68.085 ;
     RECT  98.585 67.915 98.755 68.085 ;
     RECT  102.54 67.915 102.71 68.085 ;
     RECT  105.945 67.915 106.115 68.085 ;
     RECT  106.68 67.915 106.85 68.085 ;
     RECT  112.66 67.915 112.83 68.085 ;
     RECT  113.305 67.915 113.475 68.085 ;
     RECT  117.26 67.915 117.43 68.085 ;
     RECT  15.325 68.32 15.495 68.845 ;
     RECT  42.925 68.32 43.095 68.845 ;
     RECT  70.525 68.32 70.695 68.845 ;
     RECT  98.125 68.32 98.295 68.845 ;
     RECT  29.125 72.595 29.295 73.12 ;
     RECT  56.725 72.595 56.895 73.12 ;
     RECT  84.325 72.595 84.495 73.12 ;
     RECT  111.925 72.595 112.095 73.12 ;
     RECT  1.525 73.355 1.695 73.385 ;
     RECT  29.585 73.355 29.755 73.385 ;
     RECT  10.735 73.38 10.895 73.49 ;
     RECT  28.215 73.38 28.375 73.49 ;
     RECT  58.55 73.32 58.77 73.49 ;
     RECT  60.875 73.38 61.035 73.49 ;
     RECT  62.23 73.32 62.45 73.49 ;
     RECT  81.115 73.38 81.275 73.49 ;
     RECT  112.395 73.38 112.555 73.49 ;
     RECT  1.52 73.385 1.695 73.495 ;
     RECT  19.92 73.385 20.04 73.495 ;
     RECT  29.58 73.385 29.755 73.495 ;
     RECT  61.78 73.385 61.9 73.495 ;
     RECT  65.92 73.385 66.04 73.495 ;
     RECT  71.44 73.385 71.56 73.495 ;
     RECT  78.34 73.385 78.46 73.495 ;
     RECT  97.66 73.385 97.78 73.495 ;
     RECT  111 73.385 111.12 73.495 ;
     RECT  120.66 73.385 120.78 73.495 ;
     RECT  8.915 73.38 9.025 73.5 ;
     RECT  9.375 73.38 9.485 73.5 ;
     RECT  27.775 73.38 27.885 73.5 ;
     RECT  50.775 73.38 50.885 73.5 ;
     RECT  51.695 73.38 51.805 73.5 ;
     RECT  53.515 73.39 53.675 73.5 ;
     RECT  69.635 73.38 69.745 73.5 ;
     RECT  84.815 73.38 84.925 73.5 ;
     RECT  95.855 73.38 95.965 73.5 ;
     RECT  110.115 73.38 110.225 73.5 ;
     RECT  1.525 73.495 1.695 73.525 ;
     RECT  1.985 73.355 2.155 73.525 ;
     RECT  11.46 73.355 11.63 73.525 ;
     RECT  11.645 73.355 11.815 73.525 ;
     RECT  16.06 73.355 16.23 73.525 ;
     RECT  20.385 73.355 20.555 73.525 ;
     RECT  20.845 73.355 21.015 73.525 ;
     RECT  29.585 73.495 29.755 73.525 ;
     RECT  30.04 73.355 30.21 73.525 ;
     RECT  31.7 73.355 31.87 73.525 ;
     RECT  35.565 73.355 35.735 73.525 ;
     RECT  39.52 73.355 39.69 73.525 ;
     RECT  43.385 73.355 43.555 73.525 ;
     RECT  52.86 73.355 53.03 73.525 ;
     RECT  54.7 73.355 54.87 73.525 ;
     RECT  62.245 73.49 62.415 73.525 ;
     RECT  66.66 73.355 66.83 73.525 ;
     RECT  70.985 73.355 71.155 73.525 ;
     RECT  71.905 73.355 72.075 73.525 ;
     RECT  78.805 73.355 78.975 73.525 ;
     RECT  82.03 73.355 82.2 73.525 ;
     RECT  86.625 73.355 86.795 73.525 ;
     RECT  88.465 73.355 88.635 73.525 ;
     RECT  96.56 73.355 96.73 73.525 ;
     RECT  98.86 73.355 99.03 73.525 ;
     RECT  100.425 73.355 100.595 73.525 ;
     RECT  103 73.355 103.17 73.525 ;
     RECT  107.14 73.355 107.31 73.525 ;
     RECT  111.465 73.355 111.635 73.525 ;
     RECT  113.305 73.355 113.475 73.525 ;
     RECT  57.17 73.39 57.39 73.56 ;
     RECT  15.325 73.76 15.495 74.285 ;
     RECT  42.925 73.76 43.095 74.285 ;
     RECT  70.525 73.76 70.695 74.285 ;
     RECT  98.125 73.76 98.295 74.285 ;
     RECT  29.125 78.035 29.295 78.56 ;
     RECT  56.725 78.035 56.895 78.56 ;
     RECT  84.325 78.035 84.495 78.56 ;
     RECT  111.925 78.035 112.095 78.56 ;
     RECT  83.415 78.82 83.575 78.93 ;
     RECT  119.755 78.82 119.915 78.93 ;
     RECT  1.52 78.825 1.64 78.935 ;
     RECT  7.5 78.825 7.62 78.935 ;
     RECT  29.58 78.825 29.7 78.935 ;
     RECT  57.18 78.825 57.3 78.935 ;
     RECT  70.98 78.825 71.1 78.935 ;
     RECT  94.44 78.825 94.56 78.935 ;
     RECT  97.66 78.825 97.78 78.935 ;
     RECT  111.46 78.825 111.58 78.935 ;
     RECT  120.66 78.825 120.78 78.935 ;
     RECT  5.695 78.82 5.805 78.94 ;
     RECT  33.735 78.83 33.895 78.94 ;
     RECT  1.8 78.795 1.97 78.965 ;
     RECT  1.985 78.795 2.155 78.965 ;
     RECT  7.965 78.795 8.135 78.965 ;
     RECT  9.62 78.795 9.79 78.965 ;
     RECT  13.485 78.795 13.655 78.965 ;
     RECT  15.79 78.795 15.96 78.965 ;
     RECT  19.925 78.795 20.095 78.965 ;
     RECT  21.12 78.795 21.29 78.965 ;
     RECT  24.99 78.795 25.16 78.965 ;
     RECT  29.86 78.795 30.03 78.965 ;
     RECT  30.05 78.795 30.22 78.965 ;
     RECT  31.89 78.795 32.06 78.965 ;
     RECT  34.92 78.795 35.09 78.965 ;
     RECT  39.06 78.795 39.23 78.965 ;
     RECT  42.005 78.795 42.175 78.965 ;
     RECT  43.39 78.795 43.56 78.965 ;
     RECT  47.525 78.795 47.695 78.965 ;
     RECT  49.365 78.795 49.535 78.965 ;
     RECT  55.16 78.795 55.33 78.965 ;
     RECT  57.645 78.795 57.815 78.965 ;
     RECT  59.3 78.795 59.47 78.965 ;
     RECT  63.165 78.795 63.335 78.965 ;
     RECT  67.58 78.795 67.75 78.965 ;
     RECT  71.72 78.795 71.89 78.965 ;
     RECT  75.4 78.795 75.57 78.965 ;
     RECT  75.86 78.795 76.03 78.965 ;
     RECT  79.54 78.795 79.71 78.965 ;
     RECT  79.73 78.795 79.9 78.965 ;
     RECT  84.79 78.795 84.96 78.965 ;
     RECT  87.085 78.795 87.255 78.965 ;
     RECT  89.39 78.795 89.56 78.965 ;
     RECT  93.53 78.795 93.7 78.965 ;
     RECT  94.905 78.795 95.075 78.965 ;
     RECT  98.125 78.795 98.295 78.965 ;
     RECT  98.86 78.795 99.03 78.965 ;
     RECT  102.725 78.795 102.895 78.965 ;
     RECT  105.485 78.795 105.655 78.965 ;
     RECT  107.6 78.795 107.77 78.965 ;
     RECT  112.385 78.795 112.555 78.965 ;
     RECT  113.12 78.795 113.29 78.965 ;
     RECT  117.26 78.795 117.43 78.965 ;
     RECT  71.43 78.83 71.65 79 ;
     RECT  15.325 79.2 15.495 79.725 ;
     RECT  42.925 79.2 43.095 79.725 ;
     RECT  70.525 79.2 70.695 79.725 ;
     RECT  98.125 79.2 98.295 79.725 ;
     RECT  29.125 83.475 29.295 84 ;
     RECT  56.725 83.475 56.895 84 ;
     RECT  84.325 83.475 84.495 84 ;
     RECT  111.925 83.475 112.095 84 ;
     RECT  88.935 84.26 89.095 84.37 ;
     RECT  110.555 84.26 110.715 84.37 ;
     RECT  1.52 84.265 1.64 84.375 ;
     RECT  11.18 84.265 11.3 84.375 ;
     RECT  30.5 84.265 30.62 84.375 ;
     RECT  35.1 84.265 35.22 84.375 ;
     RECT  36.94 84.265 37.06 84.375 ;
     RECT  45.22 84.265 45.34 84.375 ;
     RECT  57.18 84.265 57.3 84.375 ;
     RECT  65.92 84.265 66.04 84.375 ;
     RECT  70.06 84.265 70.18 84.375 ;
     RECT  70.98 84.265 71.1 84.375 ;
     RECT  89.84 84.265 89.96 84.375 ;
     RECT  111.46 84.265 111.58 84.375 ;
     RECT  120.66 84.265 120.78 84.375 ;
     RECT  9.375 84.26 9.485 84.38 ;
     RECT  19.035 84.26 19.145 84.38 ;
     RECT  28.695 84.26 28.805 84.38 ;
     RECT  43.415 84.26 43.525 84.38 ;
     RECT  69.155 84.27 69.315 84.38 ;
     RECT  82.955 84.27 83.115 84.38 ;
     RECT  119.755 84.27 119.915 84.38 ;
     RECT  1.8 84.235 1.97 84.405 ;
     RECT  1.985 84.235 2.155 84.405 ;
     RECT  5.665 84.235 5.835 84.405 ;
     RECT  11.645 84.235 11.815 84.405 ;
     RECT  15.785 84.235 15.955 84.405 ;
     RECT  21.12 84.235 21.29 84.405 ;
     RECT  23.42 84.235 23.59 84.405 ;
     RECT  24.985 84.235 25.155 84.405 ;
     RECT  27.29 84.235 27.46 84.405 ;
     RECT  29.585 84.235 29.755 84.405 ;
     RECT  31.24 84.235 31.41 84.405 ;
     RECT  35.565 84.235 35.735 84.405 ;
     RECT  37.68 84.235 37.85 84.405 ;
     RECT  41.55 84.235 41.72 84.405 ;
     RECT  45.685 84.235 45.855 84.405 ;
     RECT  52.59 84.235 52.76 84.405 ;
     RECT  53.045 84.235 53.215 84.405 ;
     RECT  57.645 84.235 57.815 84.405 ;
     RECT  60.405 84.235 60.575 84.405 ;
     RECT  65.01 84.235 65.18 84.405 ;
     RECT  66.385 84.235 66.555 84.405 ;
     RECT  71.445 84.235 71.615 84.405 ;
     RECT  73.745 84.235 73.915 84.405 ;
     RECT  79.08 84.235 79.25 84.405 ;
     RECT  81.105 84.235 81.275 84.405 ;
     RECT  83.87 84.235 84.04 84.405 ;
     RECT  85.06 84.235 85.23 84.405 ;
     RECT  90.31 84.235 90.48 84.405 ;
     RECT  90.77 84.235 90.94 84.405 ;
     RECT  91.685 84.235 91.855 84.405 ;
     RECT  98.585 84.235 98.755 84.405 ;
     RECT  99.045 84.235 99.215 84.405 ;
     RECT  106.68 84.235 106.85 84.405 ;
     RECT  108.245 84.235 108.415 84.405 ;
     RECT  112.66 84.235 112.83 84.405 ;
     RECT  115.88 84.235 116.05 84.405 ;
     RECT  116.8 84.235 116.97 84.405 ;
     RECT  48.89 84.27 49.11 84.44 ;
     RECT  15.325 84.64 15.495 85.165 ;
     RECT  42.925 84.64 43.095 85.165 ;
     RECT  70.525 84.64 70.695 85.165 ;
     RECT  98.125 84.64 98.295 85.165 ;
     RECT  29.125 88.915 29.295 89.44 ;
     RECT  56.725 88.915 56.895 89.44 ;
     RECT  84.325 88.915 84.495 89.44 ;
     RECT  111.925 88.915 112.095 89.44 ;
     RECT  60.405 89.675 60.575 89.705 ;
     RECT  1.52 89.705 1.64 89.71 ;
     RECT  20.855 89.7 21.015 89.81 ;
     RECT  59.035 89.7 59.195 89.81 ;
     RECT  83.415 89.7 83.575 89.81 ;
     RECT  96.755 89.7 96.915 89.81 ;
     RECT  111.015 89.7 111.175 89.81 ;
     RECT  119.755 89.7 119.915 89.81 ;
     RECT  1.52 89.71 1.695 89.815 ;
     RECT  2.44 89.705 2.56 89.815 ;
     RECT  25.9 89.705 26.02 89.815 ;
     RECT  59.94 89.705 60.06 89.815 ;
     RECT  60.4 89.705 60.575 89.815 ;
     RECT  70.06 89.705 70.18 89.815 ;
     RECT  76.04 89.705 76.16 89.815 ;
     RECT  120.66 89.705 120.78 89.815 ;
     RECT  1.535 89.815 1.695 89.82 ;
     RECT  14.415 89.71 14.575 89.82 ;
     RECT  23.175 89.7 23.285 89.82 ;
     RECT  24.995 89.71 25.155 89.82 ;
     RECT  57.215 89.7 57.325 89.82 ;
     RECT  59.495 89.71 59.655 89.82 ;
     RECT  71.935 89.7 72.045 89.82 ;
     RECT  75.135 89.71 75.295 89.82 ;
     RECT  92.155 89.71 92.315 89.82 ;
     RECT  109.195 89.7 109.305 89.82 ;
     RECT  1.985 89.675 2.155 89.845 ;
     RECT  2.905 89.675 3.075 89.845 ;
     RECT  9.345 89.675 9.515 89.845 ;
     RECT  10.54 89.675 10.71 89.845 ;
     RECT  15.79 89.675 15.96 89.845 ;
     RECT  16.98 89.675 17.15 89.845 ;
     RECT  21.765 89.675 21.935 89.845 ;
     RECT  26.365 89.675 26.535 89.845 ;
     RECT  29.585 89.675 29.755 89.845 ;
     RECT  33.73 89.675 33.9 89.845 ;
     RECT  35.565 89.675 35.735 89.845 ;
     RECT  39.52 89.675 39.69 89.845 ;
     RECT  43.385 89.675 43.555 89.845 ;
     RECT  45.5 89.675 45.67 89.845 ;
     RECT  49.37 89.675 49.54 89.845 ;
     RECT  60.405 89.815 60.575 89.845 ;
     RECT  60.865 89.675 61.035 89.845 ;
     RECT  67.77 89.675 67.94 89.845 ;
     RECT  70.99 89.675 71.16 89.845 ;
     RECT  73.745 89.675 73.915 89.845 ;
     RECT  76.505 89.675 76.675 89.845 ;
     RECT  83.87 89.675 84.04 89.845 ;
     RECT  84.785 89.675 84.955 89.845 ;
     RECT  88.005 89.675 88.175 89.845 ;
     RECT  89.39 89.675 89.56 89.845 ;
     RECT  93.07 89.675 93.24 89.845 ;
     RECT  97.665 89.675 97.835 89.845 ;
     RECT  98.585 89.675 98.755 89.845 ;
     RECT  105.3 89.675 105.47 89.845 ;
     RECT  107.785 89.675 107.955 89.845 ;
     RECT  111.465 89.675 111.635 89.845 ;
     RECT  112.385 89.675 112.555 89.845 ;
     RECT  53.03 89.71 53.25 89.88 ;
     RECT  15.325 90.08 15.495 90.605 ;
     RECT  42.925 90.08 43.095 90.605 ;
     RECT  70.525 90.08 70.695 90.605 ;
     RECT  98.125 90.08 98.295 90.605 ;
     RECT  29.125 94.355 29.295 94.88 ;
     RECT  56.725 94.355 56.895 94.88 ;
     RECT  84.325 94.355 84.495 94.88 ;
     RECT  111.925 94.355 112.095 94.88 ;
     RECT  1.555 95.14 1.665 95.145 ;
     RECT  49.36 95.145 49.48 95.15 ;
     RECT  13.495 95.14 13.655 95.25 ;
     RECT  18.555 95.14 18.715 95.25 ;
     RECT  26.835 95.14 26.995 95.25 ;
     RECT  41.095 95.14 41.255 95.25 ;
     RECT  99.055 95.14 99.215 95.25 ;
     RECT  112.395 95.14 112.555 95.25 ;
     RECT  1.52 95.145 1.665 95.255 ;
     RECT  3.36 95.145 3.48 95.255 ;
     RECT  24.52 95.145 24.64 95.255 ;
     RECT  34.18 95.145 34.3 95.255 ;
     RECT  57.18 95.145 57.3 95.255 ;
     RECT  79.72 95.145 79.84 95.255 ;
     RECT  89.84 95.145 89.96 95.255 ;
     RECT  94.44 95.145 94.56 95.255 ;
     RECT  111.46 95.145 111.58 95.255 ;
     RECT  113.3 95.145 113.42 95.255 ;
     RECT  1.555 95.255 1.665 95.26 ;
     RECT  15.815 95.14 15.925 95.26 ;
     RECT  21.795 95.14 21.905 95.26 ;
     RECT  23.615 95.15 23.775 95.26 ;
     RECT  43.395 95.15 43.555 95.26 ;
     RECT  48.455 95.15 48.615 95.26 ;
     RECT  61.355 95.14 61.465 95.26 ;
     RECT  84.815 95.14 84.925 95.26 ;
     RECT  88.035 95.14 88.145 95.26 ;
     RECT  97.215 95.15 97.375 95.26 ;
     RECT  1.985 95.115 2.155 95.285 ;
     RECT  4.1 95.115 4.27 95.285 ;
     RECT  7.965 95.115 8.135 95.285 ;
     RECT  9.62 95.115 9.79 95.285 ;
     RECT  14.68 95.115 14.85 95.285 ;
     RECT  17.9 95.115 18.07 95.285 ;
     RECT  19.465 95.115 19.635 95.285 ;
     RECT  24.99 95.115 25.16 95.285 ;
     RECT  27.74 95.115 27.91 95.285 ;
     RECT  29.59 95.115 29.76 95.285 ;
     RECT  30.505 95.115 30.675 95.285 ;
     RECT  34.65 95.115 34.82 95.285 ;
     RECT  39.7 95.115 39.875 95.285 ;
     RECT  42.005 95.115 42.175 95.285 ;
     RECT  44.58 95.115 44.75 95.285 ;
     RECT  49.825 95.115 49.995 95.285 ;
     RECT  57.46 95.115 57.63 95.285 ;
     RECT  57.645 95.115 57.815 95.285 ;
     RECT  63.165 95.115 63.335 95.285 ;
     RECT  67.58 95.115 67.75 95.285 ;
     RECT  70.985 95.115 71.155 95.285 ;
     RECT  71.45 95.115 71.62 95.285 ;
     RECT  75.86 95.115 76.03 95.285 ;
     RECT  78.62 95.115 78.79 95.285 ;
     RECT  80.19 95.115 80.36 95.285 ;
     RECT  82.485 95.115 82.655 95.285 ;
     RECT  85.705 95.115 85.875 95.285 ;
     RECT  86.63 95.115 86.8 95.285 ;
     RECT  90.58 95.115 90.75 95.285 ;
     RECT  93.34 95.115 93.51 95.285 ;
     RECT  95.18 95.115 95.35 95.285 ;
     RECT  98.585 95.115 98.755 95.285 ;
     RECT  100.24 95.115 100.41 95.285 ;
     RECT  104.105 95.115 104.275 95.285 ;
     RECT  105.945 95.115 106.115 95.285 ;
     RECT  113.765 95.115 113.935 95.285 ;
     RECT  49.35 95.15 49.57 95.32 ;
     RECT  53.03 95.15 53.25 95.32 ;
     RECT  15.325 95.52 15.495 96.045 ;
     RECT  42.925 95.52 43.095 96.045 ;
     RECT  70.525 95.52 70.695 96.045 ;
     RECT  98.125 95.52 98.295 96.045 ;
     RECT  29.125 99.795 29.295 100.32 ;
     RECT  56.725 99.795 56.895 100.32 ;
     RECT  84.325 99.795 84.495 100.32 ;
     RECT  111.925 99.795 112.095 100.32 ;
     RECT  7.515 100.58 7.675 100.69 ;
     RECT  31.435 100.58 31.595 100.69 ;
     RECT  45.695 100.58 45.855 100.69 ;
     RECT  58.575 100.58 58.735 100.69 ;
     RECT  103.655 100.58 103.815 100.69 ;
     RECT  112.395 100.58 112.555 100.69 ;
     RECT  28.2 100.585 28.32 100.695 ;
     RECT  35.56 100.585 35.68 100.695 ;
     RECT  59.48 100.585 59.6 100.695 ;
     RECT  65.92 100.585 66.04 100.695 ;
     RECT  73.28 100.585 73.4 100.695 ;
     RECT  89.84 100.585 89.96 100.695 ;
     RECT  120.66 100.585 120.78 100.695 ;
     RECT  1.555 100.58 1.665 100.7 ;
     RECT  15.795 100.59 15.955 100.7 ;
     RECT  27.315 100.58 27.425 100.7 ;
     RECT  29.615 100.58 29.725 100.7 ;
     RECT  33.275 100.59 33.435 100.7 ;
     RECT  64.115 100.58 64.225 100.7 ;
     RECT  95.395 100.58 95.505 100.7 ;
     RECT  97.215 100.59 97.375 100.7 ;
     RECT  105.955 100.59 106.115 100.7 ;
     RECT  120.215 100.59 120.375 100.7 ;
     RECT  1.8 100.555 1.97 100.725 ;
     RECT  3.64 100.555 3.81 100.725 ;
     RECT  5.665 100.555 5.835 100.725 ;
     RECT  8.425 100.555 8.595 100.725 ;
     RECT  16.705 100.555 16.875 100.725 ;
     RECT  17.625 100.555 17.795 100.725 ;
     RECT  24.34 100.555 24.51 100.725 ;
     RECT  28.67 100.555 28.84 100.725 ;
     RECT  32.345 100.555 32.515 100.725 ;
     RECT  34.19 100.555 34.36 100.725 ;
     RECT  36.025 100.555 36.195 100.725 ;
     RECT  36.935 100.555 37.105 100.725 ;
     RECT  39.705 100.555 39.875 100.725 ;
     RECT  40.17 100.555 40.34 100.725 ;
     RECT  41.54 100.555 41.71 100.725 ;
     RECT  43.385 100.555 43.555 100.725 ;
     RECT  44.31 100.555 44.48 100.725 ;
     RECT  46.6 100.555 46.77 100.725 ;
     RECT  47.985 100.555 48.155 100.725 ;
     RECT  51.21 100.555 51.38 100.725 ;
     RECT  52.13 100.555 52.3 100.725 ;
     RECT  52.86 100.555 53.03 100.725 ;
     RECT  57.19 100.555 57.36 100.725 ;
     RECT  60.22 100.555 60.39 100.725 ;
     RECT  62.245 100.555 62.415 100.725 ;
     RECT  66.385 100.555 66.555 100.725 ;
     RECT  66.66 100.555 66.83 100.725 ;
     RECT  70.99 100.555 71.16 100.725 ;
     RECT  73.745 100.555 73.915 100.725 ;
     RECT  74.665 100.555 74.835 100.725 ;
     RECT  81.38 100.555 81.55 100.725 ;
     RECT  84.785 100.555 84.955 100.725 ;
     RECT  85.25 100.555 85.42 100.725 ;
     RECT  90.31 100.555 90.48 100.725 ;
     RECT  92.145 100.555 92.315 100.725 ;
     RECT  98.585 100.555 98.755 100.725 ;
     RECT  99.78 100.555 99.95 100.725 ;
     RECT  104.565 100.555 104.735 100.725 ;
     RECT  107.14 100.555 107.31 100.725 ;
     RECT  111.005 100.555 111.175 100.725 ;
     RECT  113.305 100.555 113.475 100.725 ;
     RECT  15.325 100.96 15.495 101.485 ;
     RECT  42.925 100.96 43.095 101.485 ;
     RECT  70.525 100.96 70.695 101.485 ;
     RECT  98.125 100.96 98.295 101.485 ;
     RECT  29.125 105.235 29.295 105.76 ;
     RECT  56.725 105.235 56.895 105.76 ;
     RECT  84.325 105.235 84.495 105.76 ;
     RECT  111.925 105.235 112.095 105.76 ;
     RECT  1.525 105.995 1.695 106.025 ;
     RECT  43.39 105.995 43.56 106.025 ;
     RECT  72.825 105.995 72.995 106.025 ;
     RECT  84.785 105.995 84.955 106.025 ;
     RECT  33.735 106.02 33.895 106.13 ;
     RECT  82.955 106.02 83.115 106.13 ;
     RECT  103.195 106.02 103.355 106.13 ;
     RECT  112.395 106.02 112.555 106.13 ;
     RECT  1.52 106.025 1.695 106.135 ;
     RECT  15.78 106.025 15.9 106.135 ;
     RECT  24.06 106.025 24.18 106.135 ;
     RECT  28.66 106.025 28.78 106.135 ;
     RECT  43.38 106.025 43.56 106.135 ;
     RECT  72.82 106.025 72.995 106.135 ;
     RECT  80.18 106.025 80.3 106.135 ;
     RECT  83.86 106.025 83.98 106.135 ;
     RECT  84.78 106.025 84.955 106.135 ;
     RECT  94.44 106.025 94.56 106.135 ;
     RECT  105.48 106.025 105.6 106.135 ;
     RECT  111.46 106.025 111.58 106.135 ;
     RECT  115.14 106.025 115.26 106.135 ;
     RECT  120.66 106.025 120.78 106.135 ;
     RECT  13.515 106.02 13.625 106.14 ;
     RECT  50.755 106.03 50.915 106.14 ;
     RECT  71.015 106.02 71.125 106.14 ;
     RECT  103.675 106.02 103.785 106.14 ;
     RECT  114.235 106.03 114.395 106.14 ;
     RECT  119.755 106.03 119.915 106.14 ;
     RECT  1.525 106.135 1.695 106.165 ;
     RECT  1.985 105.995 2.155 106.165 ;
     RECT  9.62 105.995 9.79 106.165 ;
     RECT  12.565 105.995 12.735 106.165 ;
     RECT  16.25 105.995 16.42 106.165 ;
     RECT  19.93 105.995 20.1 106.165 ;
     RECT  20.39 105.995 20.56 106.165 ;
     RECT  24.525 105.995 24.7 106.165 ;
     RECT  29.86 105.995 30.03 106.165 ;
     RECT  31.89 105.995 32.06 106.165 ;
     RECT  34.65 105.995 34.82 106.165 ;
     RECT  35.565 105.995 35.735 106.165 ;
     RECT  39.705 105.995 39.875 106.165 ;
     RECT  43.39 106.135 43.56 106.165 ;
     RECT  43.845 105.995 44.015 106.165 ;
     RECT  46.15 105.995 46.32 106.165 ;
     RECT  47.985 105.995 48.155 106.165 ;
     RECT  51.665 105.995 51.835 106.165 ;
     RECT  57.19 105.995 57.36 106.165 ;
     RECT  60.41 105.995 60.58 106.165 ;
     RECT  61.785 105.995 61.955 106.165 ;
     RECT  67.31 105.995 67.48 106.165 ;
     RECT  69.14 105.995 69.31 106.165 ;
     RECT  71.44 105.995 71.61 106.165 ;
     RECT  72.825 106.135 72.995 106.165 ;
     RECT  73.285 105.995 73.455 106.165 ;
     RECT  80.65 105.995 80.82 106.165 ;
     RECT  84.785 106.135 84.955 106.165 ;
     RECT  85.25 105.995 85.42 106.165 ;
     RECT  90.58 105.995 90.75 106.165 ;
     RECT  92.42 105.995 92.59 106.165 ;
     RECT  95.18 105.995 95.35 106.165 ;
     RECT  96.29 105.995 96.46 106.165 ;
     RECT  98.59 105.995 98.76 106.165 ;
     RECT  99.32 105.995 99.49 106.165 ;
     RECT  104.105 105.995 104.275 106.165 ;
     RECT  106.22 105.995 106.39 106.165 ;
     RECT  110.36 105.995 110.53 106.165 ;
     RECT  113.305 105.995 113.475 106.165 ;
     RECT  115.88 105.995 116.05 106.165 ;
     RECT  8.87 106.03 9.09 106.2 ;
     RECT  15.325 106.4 15.495 106.925 ;
     RECT  42.925 106.4 43.095 106.925 ;
     RECT  70.525 106.4 70.695 106.925 ;
     RECT  98.125 106.4 98.295 106.925 ;
     RECT  29.125 110.675 29.295 111.2 ;
     RECT  56.725 110.675 56.895 111.2 ;
     RECT  84.325 110.675 84.495 111.2 ;
     RECT  111.925 110.675 112.095 111.2 ;
     RECT  16.715 111.46 16.875 111.57 ;
     RECT  77.435 111.46 77.595 111.57 ;
     RECT  106.875 111.46 107.035 111.57 ;
     RECT  1.52 111.465 1.64 111.575 ;
     RECT  15.78 111.465 15.9 111.575 ;
     RECT  17.62 111.465 17.74 111.575 ;
     RECT  23.6 111.465 23.72 111.575 ;
     RECT  41.08 111.465 41.2 111.575 ;
     RECT  43.38 111.465 43.5 111.575 ;
     RECT  48.9 111.465 49.02 111.575 ;
     RECT  60.4 111.465 60.52 111.575 ;
     RECT  61.78 111.465 61.9 111.575 ;
     RECT  79.26 111.465 79.38 111.575 ;
     RECT  90.76 111.465 90.88 111.575 ;
     RECT  107.78 111.465 107.9 111.575 ;
     RECT  2.915 111.47 3.075 111.58 ;
     RECT  69.615 111.47 69.775 111.58 ;
     RECT  119.315 111.46 119.425 111.58 ;
     RECT  1.985 111.435 2.155 111.605 ;
     RECT  2.445 111.435 2.615 111.605 ;
     RECT  4.1 111.435 4.27 111.605 ;
     RECT  7.965 111.435 8.135 111.605 ;
     RECT  9.345 111.435 9.515 111.605 ;
     RECT  16.245 111.435 16.415 111.605 ;
     RECT  18.09 111.435 18.26 111.605 ;
     RECT  20.85 111.435 21.02 111.605 ;
     RECT  24.065 111.435 24.235 111.605 ;
     RECT  25.26 111.435 25.43 111.605 ;
     RECT  29.585 111.435 29.755 111.605 ;
     RECT  33.725 111.435 33.895 111.605 ;
     RECT  36.945 111.435 37.115 111.605 ;
     RECT  40.63 111.435 40.8 111.605 ;
     RECT  41.55 111.435 41.72 111.605 ;
     RECT  43.845 111.435 44.015 111.605 ;
     RECT  45.225 111.435 45.395 111.605 ;
     RECT  47.065 111.435 47.235 111.605 ;
     RECT  49.79 111.435 49.96 111.605 ;
     RECT  55.81 111.435 55.98 111.605 ;
     RECT  57.185 111.435 57.36 111.605 ;
     RECT  60.87 111.435 61.04 111.605 ;
     RECT  62.25 111.435 62.42 111.605 ;
     RECT  65.465 111.435 65.635 111.605 ;
     RECT  66.385 111.435 66.555 111.605 ;
     RECT  70.985 111.435 71.155 111.605 ;
     RECT  75.125 111.435 75.295 111.605 ;
     RECT  78.35 111.435 78.52 111.605 ;
     RECT  79.725 111.435 79.895 111.605 ;
     RECT  84.79 111.435 84.96 111.605 ;
     RECT  87.085 111.435 87.255 111.605 ;
     RECT  91.225 111.435 91.395 111.605 ;
     RECT  94.445 111.435 94.615 111.605 ;
     RECT  98.585 111.435 98.755 111.605 ;
     RECT  99.505 111.435 99.675 111.605 ;
     RECT  105.945 111.435 106.115 111.605 ;
     RECT  108.245 111.435 108.415 111.605 ;
     RECT  112.39 111.435 112.56 111.605 ;
     RECT  113.305 111.435 113.475 111.605 ;
     RECT  115.42 111.435 115.59 111.605 ;
     RECT  117.26 111.435 117.43 111.605 ;
     RECT  15.325 111.84 15.495 112.365 ;
     RECT  42.925 111.84 43.095 112.365 ;
     RECT  70.525 111.84 70.695 112.365 ;
     RECT  98.125 111.84 98.295 112.365 ;
     RECT  29.125 116.115 29.295 116.64 ;
     RECT  56.725 116.115 56.895 116.64 ;
     RECT  84.325 116.115 84.495 116.64 ;
     RECT  111.925 116.115 112.095 116.64 ;
     RECT  111 116.875 111.17 116.9 ;
     RECT  112.38 116.905 112.5 116.91 ;
     RECT  7.515 116.9 7.675 117.01 ;
     RECT  18.095 116.9 18.255 117.01 ;
     RECT  26.375 116.9 26.535 117.01 ;
     RECT  111 116.9 111.175 117.01 ;
     RECT  120.215 116.9 120.375 117.01 ;
     RECT  1.52 116.905 1.64 117.015 ;
     RECT  2.9 116.905 3.02 117.015 ;
     RECT  15.78 116.905 15.9 117.015 ;
     RECT  24.52 116.905 24.64 117.015 ;
     RECT  27.28 116.905 27.4 117.015 ;
     RECT  29.12 116.905 29.24 117.015 ;
     RECT  41.54 116.905 41.66 117.015 ;
     RECT  68.22 116.905 68.34 117.015 ;
     RECT  70.06 116.905 70.18 117.015 ;
     RECT  72.36 116.905 72.48 117.015 ;
     RECT  112.38 116.91 112.555 117.015 ;
     RECT  113.3 116.905 113.42 117.015 ;
     RECT  9.375 116.9 9.485 117.02 ;
     RECT  41.115 116.9 41.225 117.02 ;
     RECT  112.395 117.015 112.555 117.02 ;
     RECT  1.985 116.875 2.155 117.045 ;
     RECT  2.445 116.875 2.615 117.045 ;
     RECT  3.64 116.875 3.81 117.045 ;
     RECT  8.425 116.875 8.595 117.045 ;
     RECT  11.46 116.875 11.63 117.045 ;
     RECT  16.52 116.875 16.69 117.045 ;
     RECT  19.005 116.875 19.175 117.045 ;
     RECT  20.66 116.875 20.83 117.045 ;
     RECT  24.99 116.875 25.16 117.045 ;
     RECT  27.74 116.875 27.91 117.045 ;
     RECT  29.59 116.875 29.76 117.045 ;
     RECT  29.86 116.875 30.03 117.045 ;
     RECT  33.73 116.875 33.9 117.045 ;
     RECT  34.185 116.875 34.355 117.045 ;
     RECT  37.87 116.875 38.04 117.045 ;
     RECT  42.01 116.875 42.18 117.045 ;
     RECT  43.385 116.875 43.56 117.045 ;
     RECT  46.605 116.875 46.775 117.045 ;
     RECT  47.525 116.875 47.695 117.045 ;
     RECT  49.83 116.875 50 117.045 ;
     RECT  50.74 116.875 50.91 117.045 ;
     RECT  52.125 116.875 52.295 117.045 ;
     RECT  53.045 116.875 53.215 117.045 ;
     RECT  57.185 116.875 57.355 117.045 ;
     RECT  60.865 116.875 61.04 117.045 ;
     RECT  65.465 116.875 65.635 117.045 ;
     RECT  68.69 116.875 68.86 117.045 ;
     RECT  70.99 116.875 71.16 117.045 ;
     RECT  72.83 116.875 73 117.045 ;
     RECT  73.75 116.875 73.92 117.045 ;
     RECT  80.185 116.875 80.355 117.045 ;
     RECT  81.105 116.875 81.275 117.045 ;
     RECT  84.785 116.875 84.955 117.045 ;
     RECT  89.39 116.875 89.56 117.045 ;
     RECT  92.145 116.875 92.315 117.045 ;
     RECT  93.99 116.875 94.16 117.045 ;
     RECT  98.86 116.875 99.03 117.045 ;
     RECT  99.505 116.875 99.675 117.045 ;
     RECT  103 116.875 103.17 117.045 ;
     RECT  107.14 116.875 107.31 117.045 ;
     RECT  111 117.01 111.17 117.045 ;
     RECT  112.845 116.875 113.015 117.045 ;
     RECT  113.765 116.875 113.935 117.045 ;
     RECT  15.325 117.28 15.495 117.805 ;
     RECT  42.925 117.28 43.095 117.805 ;
     RECT  70.525 117.28 70.695 117.805 ;
     RECT  98.125 117.28 98.295 117.805 ;
     RECT  29.125 121.555 29.295 122.08 ;
     RECT  56.725 121.555 56.895 122.08 ;
     RECT  84.325 121.555 84.495 122.08 ;
     RECT  111.925 121.555 112.095 122.08 ;
     RECT  17.175 122.34 17.335 122.45 ;
     RECT  28.215 122.34 28.375 122.45 ;
     RECT  29.595 122.34 29.755 122.45 ;
     RECT  43.855 122.34 44.015 122.45 ;
     RECT  67.775 122.34 67.935 122.45 ;
     RECT  112.395 122.34 112.555 122.45 ;
     RECT  1.52 122.345 1.64 122.455 ;
     RECT  25.9 122.345 26.02 122.455 ;
     RECT  30.5 122.345 30.62 122.455 ;
     RECT  35.1 122.345 35.22 122.455 ;
     RECT  53.5 122.345 53.62 122.455 ;
     RECT  56.26 122.345 56.38 122.455 ;
     RECT  70.98 122.345 71.1 122.455 ;
     RECT  76.5 122.345 76.62 122.455 ;
     RECT  104.1 122.345 104.22 122.455 ;
     RECT  120.66 122.345 120.78 122.455 ;
     RECT  9.375 122.34 9.485 122.46 ;
     RECT  23.175 122.34 23.285 122.46 ;
     RECT  24.995 122.35 25.155 122.46 ;
     RECT  45.695 122.35 45.855 122.46 ;
     RECT  119.315 122.34 119.425 122.46 ;
     RECT  1.985 122.315 2.155 122.485 ;
     RECT  9.62 122.315 9.79 122.485 ;
     RECT  11.46 122.315 11.63 122.485 ;
     RECT  15.785 122.315 15.955 122.485 ;
     RECT  18.36 122.315 18.53 122.485 ;
     RECT  22.5 122.315 22.67 122.485 ;
     RECT  26.365 122.315 26.535 122.485 ;
     RECT  30.96 122.315 31.13 122.485 ;
     RECT  33.265 122.315 33.435 122.485 ;
     RECT  33.72 122.315 33.89 122.485 ;
     RECT  34.18 122.315 34.35 122.485 ;
     RECT  35.565 122.315 35.735 122.485 ;
     RECT  36.485 122.315 36.655 122.485 ;
     RECT  43.39 122.315 43.56 122.485 ;
     RECT  44.765 122.315 44.935 122.485 ;
     RECT  46.605 122.315 46.775 122.485 ;
     RECT  53.97 122.315 54.14 122.485 ;
     RECT  55.805 122.315 55.975 122.485 ;
     RECT  57.19 122.315 57.36 122.485 ;
     RECT  58.565 122.315 58.735 122.485 ;
     RECT  59.49 122.315 59.66 122.485 ;
     RECT  61.785 122.315 61.955 122.485 ;
     RECT  68.685 122.315 68.855 122.485 ;
     RECT  71.45 122.315 71.62 122.485 ;
     RECT  73.285 122.315 73.455 122.485 ;
     RECT  76.965 122.315 77.135 122.485 ;
     RECT  78.62 122.315 78.79 122.485 ;
     RECT  82.485 122.315 82.655 122.485 ;
     RECT  84.785 122.315 84.955 122.485 ;
     RECT  89.85 122.315 90.02 122.485 ;
     RECT  92.15 122.315 92.32 122.485 ;
     RECT  94.26 122.315 94.43 122.485 ;
     RECT  96.75 122.315 96.92 122.485 ;
     RECT  98.585 122.315 98.76 122.485 ;
     RECT  102.265 122.315 102.435 122.485 ;
     RECT  103.65 122.315 103.82 122.485 ;
     RECT  104.565 122.315 104.735 122.485 ;
     RECT  108.245 122.315 108.415 122.485 ;
     RECT  111.925 122.315 112.095 122.485 ;
     RECT  113.305 122.315 113.475 122.485 ;
     RECT  13.47 122.35 13.69 122.52 ;
     RECT  15.325 122.72 15.495 123.245 ;
     RECT  42.925 122.72 43.095 123.245 ;
     RECT  70.525 122.72 70.695 123.245 ;
     RECT  98.125 122.72 98.295 123.245 ;
     RECT  29.125 126.995 29.295 127.52 ;
     RECT  56.725 126.995 56.895 127.52 ;
     RECT  84.325 126.995 84.495 127.52 ;
     RECT  111.925 126.995 112.095 127.52 ;
     RECT  1.52 127.785 1.64 127.79 ;
     RECT  45.23 127.755 45.4 127.79 ;
     RECT  36.955 127.78 37.115 127.89 ;
     RECT  66.395 127.78 66.555 127.89 ;
     RECT  81.575 127.78 81.735 127.89 ;
     RECT  1.52 127.79 1.695 127.895 ;
     RECT  9.34 127.785 9.46 127.895 ;
     RECT  21.3 127.785 21.42 127.895 ;
     RECT  48.9 127.785 49.02 127.895 ;
     RECT  57.18 127.785 57.3 127.895 ;
     RECT  74.66 127.785 74.78 127.895 ;
     RECT  77.88 127.785 78 127.895 ;
     RECT  84.78 127.785 84.9 127.895 ;
     RECT  89.38 127.785 89.5 127.895 ;
     RECT  105.02 127.785 105.14 127.895 ;
     RECT  109.62 127.785 109.74 127.895 ;
     RECT  115.14 127.785 115.26 127.895 ;
     RECT  120.66 127.785 120.78 127.895 ;
     RECT  1.535 127.895 1.695 127.9 ;
     RECT  15.795 127.79 15.955 127.9 ;
     RECT  43.415 127.78 43.525 127.9 ;
     RECT  69.615 127.79 69.775 127.9 ;
     RECT  97.215 127.79 97.375 127.9 ;
     RECT  114.235 127.79 114.395 127.9 ;
     RECT  119.755 127.79 119.915 127.9 ;
     RECT  1.985 127.755 2.155 127.925 ;
     RECT  2.72 127.755 2.89 127.925 ;
     RECT  6.585 127.755 6.755 127.925 ;
     RECT  9.805 127.755 9.975 127.925 ;
     RECT  14.865 127.755 15.035 127.925 ;
     RECT  16.705 127.755 16.875 127.925 ;
     RECT  17.44 127.755 17.61 127.925 ;
     RECT  21.765 127.755 21.935 127.925 ;
     RECT  24.065 127.755 24.235 127.925 ;
     RECT  29.86 127.755 30.03 127.925 ;
     RECT  33.725 127.755 33.895 127.925 ;
     RECT  34.64 127.755 34.81 127.925 ;
     RECT  37.865 127.755 38.035 127.925 ;
     RECT  41.09 127.755 41.26 127.925 ;
     RECT  49.365 127.755 49.535 127.925 ;
     RECT  52.86 127.755 53.03 127.925 ;
     RECT  56.725 127.755 56.895 127.925 ;
     RECT  57.645 127.755 57.815 127.925 ;
     RECT  65.47 127.755 65.64 127.925 ;
     RECT  67.31 127.755 67.48 127.925 ;
     RECT  70.99 127.755 71.16 127.925 ;
     RECT  75.13 127.755 75.3 127.925 ;
     RECT  78.345 127.755 78.515 127.925 ;
     RECT  82.485 127.755 82.655 127.925 ;
     RECT  85.25 127.755 85.42 127.925 ;
     RECT  85.705 127.755 85.875 127.925 ;
     RECT  89.85 127.755 90.02 127.925 ;
     RECT  93.07 127.755 93.24 127.925 ;
     RECT  97.665 127.755 97.835 127.925 ;
     RECT  98.585 127.755 98.755 127.925 ;
     RECT  105.49 127.755 105.66 127.925 ;
     RECT  105.945 127.755 106.115 127.925 ;
     RECT  108.245 127.755 108.415 127.925 ;
     RECT  110.36 127.755 110.53 127.925 ;
     RECT  112.66 127.755 112.83 127.925 ;
     RECT  115.88 127.755 116.05 127.925 ;
     RECT  116.8 127.755 116.97 127.925 ;
     RECT  45.21 127.79 45.43 127.96 ;
     RECT  15.325 128.16 15.495 128.685 ;
     RECT  42.925 128.16 43.095 128.685 ;
     RECT  70.525 128.16 70.695 128.685 ;
     RECT  98.125 128.16 98.295 128.685 ;
     RECT  29.125 132.435 29.295 132.96 ;
     RECT  56.725 132.435 56.895 132.96 ;
     RECT  84.325 132.435 84.495 132.96 ;
     RECT  111.925 132.435 112.095 132.96 ;
     RECT  18.555 133.22 18.715 133.33 ;
     RECT  100.435 133.22 100.595 133.33 ;
     RECT  112.395 133.22 112.555 133.33 ;
     RECT  2.44 133.225 2.56 133.335 ;
     RECT  4.28 133.225 4.4 133.335 ;
     RECT  10.72 133.225 10.84 133.335 ;
     RECT  17.62 133.225 17.74 133.335 ;
     RECT  19.46 133.225 19.58 133.335 ;
     RECT  29.58 133.225 29.7 133.335 ;
     RECT  45.68 133.225 45.8 133.335 ;
     RECT  56.26 133.225 56.38 133.335 ;
     RECT  56.72 133.225 56.84 133.335 ;
     RECT  63.16 133.225 63.28 133.335 ;
     RECT  98.58 133.225 98.7 133.335 ;
     RECT  103.18 133.225 103.3 133.335 ;
     RECT  111.46 133.225 111.58 133.335 ;
     RECT  112.84 133.225 112.96 133.335 ;
     RECT  120.66 133.225 120.78 133.335 ;
     RECT  15.815 133.22 15.925 133.34 ;
     RECT  34.655 133.23 34.815 133.34 ;
     RECT  42.955 133.22 43.065 133.34 ;
     RECT  55.815 133.23 55.975 133.34 ;
     RECT  61.355 133.22 61.465 133.34 ;
     RECT  69.615 133.23 69.775 133.34 ;
     RECT  79.295 133.22 79.405 133.34 ;
     RECT  86.195 133.22 86.305 133.34 ;
     RECT  95.375 133.23 95.535 133.34 ;
     RECT  109.655 133.22 109.765 133.34 ;
     RECT  111.035 133.22 111.145 133.34 ;
     RECT  1.525 133.195 1.695 133.365 ;
     RECT  3.825 133.195 3.995 133.365 ;
     RECT  5.02 133.195 5.19 133.365 ;
     RECT  8.885 133.195 9.055 133.365 ;
     RECT  11.46 133.195 11.63 133.365 ;
     RECT  18.36 133.195 18.53 133.365 ;
     RECT  19.925 133.195 20.095 133.365 ;
     RECT  22.225 133.195 22.395 133.365 ;
     RECT  27.29 133.195 27.46 133.365 ;
     RECT  30.04 133.195 30.21 133.365 ;
     RECT  31.7 133.195 31.87 133.365 ;
     RECT  31.89 133.195 32.06 133.365 ;
     RECT  35.565 133.195 35.735 133.365 ;
     RECT  43.38 133.195 43.55 133.365 ;
     RECT  44.77 133.195 44.94 133.365 ;
     RECT  46.145 133.195 46.315 133.365 ;
     RECT  48.905 133.195 49.075 133.365 ;
     RECT  57.19 133.195 57.36 133.365 ;
     RECT  63.63 133.195 63.8 133.365 ;
     RECT  65.005 133.195 65.175 133.365 ;
     RECT  66.39 133.195 66.56 133.365 ;
     RECT  71.26 133.195 71.43 133.365 ;
     RECT  72.83 133.195 73 133.365 ;
     RECT  75.4 133.195 75.57 133.365 ;
     RECT  80.46 133.195 80.63 133.365 ;
     RECT  81.11 133.195 81.28 133.365 ;
     RECT  84.785 133.195 84.955 133.365 ;
     RECT  86.9 133.195 87.07 133.365 ;
     RECT  88.01 133.195 88.18 133.365 ;
     RECT  90.77 133.195 90.94 133.365 ;
     RECT  92.14 133.195 92.31 133.365 ;
     RECT  93.53 133.195 93.7 133.365 ;
     RECT  94.91 133.195 95.08 133.365 ;
     RECT  96.29 133.195 96.46 133.365 ;
     RECT  99.04 133.195 99.21 133.365 ;
     RECT  99.32 133.195 99.49 133.365 ;
     RECT  101.62 133.195 101.79 133.365 ;
     RECT  103.645 133.195 103.815 133.365 ;
     RECT  105.76 133.195 105.93 133.365 ;
     RECT  113.305 133.195 113.475 133.365 ;
     RECT  15.325 133.6 15.495 134.125 ;
     RECT  42.925 133.6 43.095 134.125 ;
     RECT  70.525 133.6 70.695 134.125 ;
     RECT  98.125 133.6 98.295 134.125 ;
     RECT  29.125 137.875 29.295 138.4 ;
     RECT  56.725 137.875 56.895 138.4 ;
     RECT  84.325 137.875 84.495 138.4 ;
     RECT  111.925 137.875 112.095 138.4 ;
     RECT  70.065 138.635 70.235 138.665 ;
     RECT  88.495 138.66 88.605 138.665 ;
     RECT  55.355 138.66 55.515 138.77 ;
     RECT  68.695 138.66 68.855 138.77 ;
     RECT  81.575 138.66 81.735 138.77 ;
     RECT  1.52 138.665 1.64 138.775 ;
     RECT  9.34 138.665 9.46 138.775 ;
     RECT  15.78 138.665 15.9 138.775 ;
     RECT  24.52 138.665 24.64 138.775 ;
     RECT  44.3 138.665 44.42 138.775 ;
     RECT  45.68 138.665 45.8 138.775 ;
     RECT  56.26 138.665 56.38 138.775 ;
     RECT  69.6 138.665 69.72 138.775 ;
     RECT  70.06 138.665 70.235 138.775 ;
     RECT  88.46 138.665 88.605 138.775 ;
     RECT  90.3 138.665 90.42 138.775 ;
     RECT  97.66 138.665 97.78 138.775 ;
     RECT  98.58 138.665 98.7 138.775 ;
     RECT  102.72 138.665 102.84 138.775 ;
     RECT  104.1 138.665 104.22 138.775 ;
     RECT  116.06 138.665 116.18 138.775 ;
     RECT  120.66 138.665 120.78 138.775 ;
     RECT  2.915 138.67 3.075 138.78 ;
     RECT  29.615 138.66 29.725 138.78 ;
     RECT  42.015 138.67 42.175 138.78 ;
     RECT  42.955 138.66 43.065 138.78 ;
     RECT  43.395 138.67 43.555 138.78 ;
     RECT  53.535 138.66 53.645 138.78 ;
     RECT  69.155 138.67 69.315 138.78 ;
     RECT  88.495 138.775 88.605 138.78 ;
     RECT  1.985 138.635 2.155 138.805 ;
     RECT  2.445 138.635 2.615 138.805 ;
     RECT  4.1 138.635 4.27 138.805 ;
     RECT  7.965 138.635 8.135 138.805 ;
     RECT  9.805 138.635 9.975 138.805 ;
     RECT  16.25 138.635 16.42 138.805 ;
     RECT  17.165 138.635 17.335 138.805 ;
     RECT  19.005 138.635 19.175 138.805 ;
     RECT  25.26 138.635 25.43 138.805 ;
     RECT  28.205 138.635 28.375 138.805 ;
     RECT  30.51 138.635 30.68 138.805 ;
     RECT  31.7 138.635 31.87 138.805 ;
     RECT  34.65 138.635 34.82 138.805 ;
     RECT  35.565 138.635 35.735 138.805 ;
     RECT  44.765 138.635 44.935 138.805 ;
     RECT  46.145 138.635 46.315 138.805 ;
     RECT  52.125 138.635 52.295 138.805 ;
     RECT  57.185 138.635 57.355 138.805 ;
     RECT  59.485 138.635 59.655 138.805 ;
     RECT  64.82 138.635 64.99 138.805 ;
     RECT  70.065 138.775 70.235 138.805 ;
     RECT  70.985 138.635 71.155 138.805 ;
     RECT  77.43 138.635 77.6 138.805 ;
     RECT  78.62 138.635 78.79 138.805 ;
     RECT  82.485 138.635 82.655 138.805 ;
     RECT  84.6 138.635 84.77 138.805 ;
     RECT  84.785 138.635 84.955 138.805 ;
     RECT  88.925 138.635 89.095 138.805 ;
     RECT  91.04 138.635 91.21 138.805 ;
     RECT  94.905 138.635 95.075 138.805 ;
     RECT  96.28 138.635 96.45 138.805 ;
     RECT  98.86 138.635 99.03 138.805 ;
     RECT  99.04 138.635 99.21 138.805 ;
     RECT  103.19 138.635 103.36 138.805 ;
     RECT  104.565 138.635 104.735 138.805 ;
     RECT  107.785 138.635 107.955 138.805 ;
     RECT  112.385 138.635 112.555 138.805 ;
     RECT  116.8 138.635 116.97 138.805 ;
     RECT  116.985 138.635 117.155 138.805 ;
     RECT  100.41 138.67 100.63 138.84 ;
     RECT  15.325 139.04 15.495 139.565 ;
     RECT  42.925 139.04 43.095 139.565 ;
     RECT  70.525 139.04 70.695 139.565 ;
     RECT  98.125 139.04 98.295 139.565 ;
     RECT  29.125 143.315 29.295 143.84 ;
     RECT  56.725 143.315 56.895 143.84 ;
     RECT  84.325 143.315 84.495 143.84 ;
     RECT  111.925 143.315 112.095 143.84 ;
     RECT  88.92 144.075 89.09 144.11 ;
     RECT  15.335 144.1 15.495 144.21 ;
     RECT  51.215 144.1 51.375 144.21 ;
     RECT  111.015 144.1 111.175 144.21 ;
     RECT  18.54 144.105 18.66 144.215 ;
     RECT  25.9 144.105 26.02 144.215 ;
     RECT  52.12 144.105 52.24 144.215 ;
     RECT  62.7 144.105 62.82 144.215 ;
     RECT  76.5 144.105 76.62 144.215 ;
     RECT  120.66 144.105 120.78 144.215 ;
     RECT  14.415 144.11 14.575 144.22 ;
     RECT  15.815 144.1 15.925 144.22 ;
     RECT  17.635 144.11 17.795 144.22 ;
     RECT  43.395 144.11 43.555 144.22 ;
     RECT  49.395 144.1 49.505 144.22 ;
     RECT  55.835 144.1 55.945 144.22 ;
     RECT  57.215 144.1 57.325 144.22 ;
     RECT  61.795 144.11 61.955 144.22 ;
     RECT  75.155 144.1 75.265 144.22 ;
     RECT  88.92 144.11 89.095 144.22 ;
     RECT  1.525 144.075 1.695 144.245 ;
     RECT  2.445 144.075 2.615 144.245 ;
     RECT  3.18 144.075 3.35 144.245 ;
     RECT  7.045 144.075 7.215 144.245 ;
     RECT  11.46 144.075 11.63 144.245 ;
     RECT  16.245 144.075 16.415 144.245 ;
     RECT  19.005 144.075 19.175 144.245 ;
     RECT  26.37 144.075 26.54 144.245 ;
     RECT  28.205 144.075 28.375 144.245 ;
     RECT  29.59 144.075 29.76 144.245 ;
     RECT  34.65 144.075 34.82 144.245 ;
     RECT  35.565 144.075 35.735 144.245 ;
     RECT  42.005 144.075 42.175 144.245 ;
     RECT  44.305 144.075 44.475 144.245 ;
     RECT  51.94 144.075 52.11 144.245 ;
     RECT  52.86 144.075 53.03 144.245 ;
     RECT  57.65 144.075 57.82 144.245 ;
     RECT  59.025 144.075 59.195 144.245 ;
     RECT  63.165 144.075 63.335 144.245 ;
     RECT  66.39 144.075 66.56 144.245 ;
     RECT  70.99 144.075 71.16 144.245 ;
     RECT  76.965 144.075 77.135 144.245 ;
     RECT  77.885 144.075 78.055 144.245 ;
     RECT  85.06 144.075 85.23 144.245 ;
     RECT  85.245 144.075 85.415 144.245 ;
     RECT  88.92 144.22 89.09 144.245 ;
     RECT  89.85 144.075 90.02 144.245 ;
     RECT  90.305 144.075 90.475 144.245 ;
     RECT  92.88 144.075 93.05 144.245 ;
     RECT  96.74 144.075 96.91 144.245 ;
     RECT  97.665 144.075 97.835 144.245 ;
     RECT  98.585 144.075 98.755 144.245 ;
     RECT  105.03 144.075 105.2 144.245 ;
     RECT  105.94 144.075 106.11 144.245 ;
     RECT  107.14 144.075 107.31 144.245 ;
     RECT  107.6 144.075 107.77 144.245 ;
     RECT  111.47 144.075 111.64 144.245 ;
     RECT  112.66 144.075 112.83 144.245 ;
     RECT  113.305 144.075 113.475 144.245 ;
     RECT  116.8 144.075 116.97 144.245 ;
     RECT  15.325 144.48 15.495 145.005 ;
     RECT  42.925 144.48 43.095 145.005 ;
     RECT  70.525 144.48 70.695 145.005 ;
     RECT  98.125 144.48 98.295 145.005 ;
     RECT  29.125 148.755 29.295 149.28 ;
     RECT  56.725 148.755 56.895 149.28 ;
     RECT  84.325 148.755 84.495 149.28 ;
     RECT  111.925 148.755 112.095 149.28 ;
     RECT  54.915 149.54 55.025 149.545 ;
     RECT  70.065 149.515 70.235 149.545 ;
     RECT  46.615 149.54 46.775 149.65 ;
     RECT  69.155 149.54 69.315 149.65 ;
     RECT  83.415 149.54 83.575 149.65 ;
     RECT  99.055 149.54 99.215 149.65 ;
     RECT  13.94 149.545 14.06 149.655 ;
     RECT  14.86 149.545 14.98 149.655 ;
     RECT  18.54 149.545 18.66 149.655 ;
     RECT  33.72 149.545 33.84 149.655 ;
     RECT  42.46 149.545 42.58 149.655 ;
     RECT  54.88 149.545 55.025 149.655 ;
     RECT  57.18 149.545 57.3 149.655 ;
     RECT  65.46 149.545 65.58 149.655 ;
     RECT  70.06 149.545 70.235 149.655 ;
     RECT  79.26 149.545 79.38 149.655 ;
     RECT  104.1 149.545 104.22 149.655 ;
     RECT  116.06 149.545 116.18 149.655 ;
     RECT  120.66 149.545 120.78 149.655 ;
     RECT  1.555 149.54 1.665 149.66 ;
     RECT  12.135 149.54 12.245 149.66 ;
     RECT  15.815 149.54 15.925 149.66 ;
     RECT  17.635 149.55 17.795 149.66 ;
     RECT  41.555 149.55 41.715 149.66 ;
     RECT  54.915 149.655 55.025 149.66 ;
     RECT  62.735 149.54 62.845 149.66 ;
     RECT  64.555 149.55 64.715 149.66 ;
     RECT  77.455 149.54 77.565 149.66 ;
     RECT  120.215 149.55 120.375 149.66 ;
     RECT  3.365 149.515 3.535 149.685 ;
     RECT  4.285 149.515 4.455 149.685 ;
     RECT  11.645 149.515 11.815 149.685 ;
     RECT  14.405 149.515 14.575 149.685 ;
     RECT  19.005 149.515 19.175 149.685 ;
     RECT  21.765 149.515 21.935 149.685 ;
     RECT  26.365 149.515 26.535 149.685 ;
     RECT  29.58 149.515 29.75 149.685 ;
     RECT  31.885 149.515 32.055 149.685 ;
     RECT  34.185 149.515 34.355 149.685 ;
     RECT  39.245 149.515 39.415 149.685 ;
     RECT  43.39 149.515 43.56 149.685 ;
     RECT  45.225 149.515 45.395 149.685 ;
     RECT  47.525 149.515 47.695 149.685 ;
     RECT  55.345 149.515 55.515 149.685 ;
     RECT  57.645 149.515 57.815 149.685 ;
     RECT  65.01 149.515 65.18 149.685 ;
     RECT  66.2 149.515 66.37 149.685 ;
     RECT  70.065 149.655 70.235 149.685 ;
     RECT  70.985 149.515 71.155 149.685 ;
     RECT  78.62 149.515 78.79 149.685 ;
     RECT  79.725 149.515 79.895 149.685 ;
     RECT  82.76 149.515 82.93 149.685 ;
     RECT  84.79 149.515 84.96 149.685 ;
     RECT  86.63 149.515 86.8 149.685 ;
     RECT  89.385 149.515 89.555 149.685 ;
     RECT  91.23 149.515 91.4 149.685 ;
     RECT  94.445 149.515 94.615 149.685 ;
     RECT  98.59 149.515 98.76 149.685 ;
     RECT  100.24 149.515 100.41 149.685 ;
     RECT  103.19 149.515 103.36 149.685 ;
     RECT  104.565 149.515 104.735 149.685 ;
     RECT  105.025 149.515 105.195 149.685 ;
     RECT  112.385 149.515 112.555 149.685 ;
     RECT  113.305 149.515 113.475 149.685 ;
     RECT  116.525 149.515 116.695 149.685 ;
     RECT  15.325 149.92 15.495 150.445 ;
     RECT  42.925 149.92 43.095 150.445 ;
     RECT  70.525 149.92 70.695 150.445 ;
     RECT  98.125 149.92 98.295 150.445 ;
     RECT  29.125 154.195 29.295 154.72 ;
     RECT  56.725 154.195 56.895 154.72 ;
     RECT  84.325 154.195 84.495 154.72 ;
     RECT  111.925 154.195 112.095 154.72 ;
     RECT  70.065 154.955 70.235 154.985 ;
     RECT  1.555 154.98 1.665 154.99 ;
     RECT  18.555 154.98 18.715 155.09 ;
     RECT  81.115 154.98 81.275 155.09 ;
     RECT  91.235 154.98 91.395 155.09 ;
     RECT  2.44 154.985 2.56 155.095 ;
     RECT  3.36 154.985 3.48 155.095 ;
     RECT  38.32 154.985 38.44 155.095 ;
     RECT  55.8 154.985 55.92 155.095 ;
     RECT  56.26 154.985 56.38 155.095 ;
     RECT  70.06 154.985 70.235 155.095 ;
     RECT  71.9 154.985 72.02 155.095 ;
     RECT  76.5 154.985 76.62 155.095 ;
     RECT  82.02 154.985 82.14 155.095 ;
     RECT  88.92 154.985 89.04 155.095 ;
     RECT  99.5 154.985 99.62 155.095 ;
     RECT  108.7 154.985 108.82 155.095 ;
     RECT  112.38 154.985 112.5 155.095 ;
     RECT  120.66 154.985 120.78 155.095 ;
     RECT  1.535 154.99 1.695 155.1 ;
     RECT  15.815 154.98 15.925 155.1 ;
     RECT  21.775 154.99 21.935 155.1 ;
     RECT  29.615 154.98 29.725 155.1 ;
     RECT  37.415 154.99 37.575 155.1 ;
     RECT  43.395 154.99 43.555 155.1 ;
     RECT  70.995 154.99 71.155 155.1 ;
     RECT  98.595 154.99 98.755 155.1 ;
     RECT  3.18 154.955 3.35 155.125 ;
     RECT  3.825 154.955 3.995 155.125 ;
     RECT  7.32 154.955 7.49 155.125 ;
     RECT  11.185 154.955 11.355 155.125 ;
     RECT  11.46 154.955 11.63 155.125 ;
     RECT  17.9 154.955 18.07 155.125 ;
     RECT  19.465 154.955 19.635 155.125 ;
     RECT  22.685 154.955 22.855 155.125 ;
     RECT  26.82 154.955 26.99 155.125 ;
     RECT  30.045 154.955 30.215 155.125 ;
     RECT  31.7 154.955 31.87 155.125 ;
     RECT  35.565 154.955 35.735 155.125 ;
     RECT  39.06 154.955 39.23 155.125 ;
     RECT  44.58 154.955 44.75 155.125 ;
     RECT  44.765 154.955 44.935 155.125 ;
     RECT  48.445 154.955 48.615 155.125 ;
     RECT  48.72 154.955 48.89 155.125 ;
     RECT  56.54 154.955 56.71 155.125 ;
     RECT  60.405 154.955 60.575 155.125 ;
     RECT  60.865 154.955 61.035 155.125 ;
     RECT  70.065 155.095 70.235 155.125 ;
     RECT  72.64 154.955 72.81 155.125 ;
     RECT  76.965 154.955 77.135 155.125 ;
     RECT  77.425 154.955 77.595 155.125 ;
     RECT  82.485 154.955 82.655 155.125 ;
     RECT  84.325 154.955 84.495 155.125 ;
     RECT  85.06 154.955 85.23 155.125 ;
     RECT  88.01 154.955 88.18 155.125 ;
     RECT  89.39 154.955 89.56 155.125 ;
     RECT  90.765 154.955 90.935 155.125 ;
     RECT  92.145 154.955 92.315 155.125 ;
     RECT  99.965 154.955 100.135 155.125 ;
     RECT  101.345 154.955 101.515 155.125 ;
     RECT  103.92 154.955 104.09 155.125 ;
     RECT  108.06 154.955 108.23 155.125 ;
     RECT  109.17 154.955 109.34 155.125 ;
     RECT  111.93 154.955 112.1 155.125 ;
     RECT  112.845 154.955 113.015 155.125 ;
     RECT  116.8 154.955 116.97 155.125 ;
     RECT  116.985 154.955 117.155 155.125 ;
     RECT  52.57 154.99 52.79 155.16 ;
     RECT  57.17 154.99 57.39 155.16 ;
     RECT  15.325 155.36 15.495 155.885 ;
     RECT  42.925 155.36 43.095 155.885 ;
     RECT  70.525 155.36 70.695 155.885 ;
     RECT  98.125 155.36 98.295 155.885 ;
     RECT  29.125 159.635 29.295 160.16 ;
     RECT  56.725 159.635 56.895 160.16 ;
     RECT  84.325 159.635 84.495 160.16 ;
     RECT  111.925 159.635 112.095 160.16 ;
     RECT  1.535 160.42 1.695 160.425 ;
     RECT  111.465 160.395 111.635 160.425 ;
     RECT  1.52 160.425 1.695 160.53 ;
     RECT  27.755 160.42 27.915 160.53 ;
     RECT  29.595 160.42 29.755 160.53 ;
     RECT  66.37 160.36 66.59 160.53 ;
     RECT  96.755 160.42 96.915 160.53 ;
     RECT  105.495 160.42 105.655 160.53 ;
     RECT  110.555 160.42 110.715 160.53 ;
     RECT  112.395 160.42 112.555 160.53 ;
     RECT  1.52 160.53 1.64 160.535 ;
     RECT  28.66 160.425 28.78 160.535 ;
     RECT  40.16 160.425 40.28 160.535 ;
     RECT  61.78 160.425 61.9 160.535 ;
     RECT  70.06 160.425 70.18 160.535 ;
     RECT  82.48 160.425 82.6 160.535 ;
     RECT  97.66 160.425 97.78 160.535 ;
     RECT  99.5 160.425 99.62 160.535 ;
     RECT  111.46 160.425 111.635 160.535 ;
     RECT  120.66 160.425 120.78 160.535 ;
     RECT  9.375 160.42 9.485 160.54 ;
     RECT  25.935 160.42 26.045 160.54 ;
     RECT  32.835 160.42 32.945 160.54 ;
     RECT  34.655 160.43 34.815 160.54 ;
     RECT  59.055 160.42 59.165 160.54 ;
     RECT  60.875 160.43 61.035 160.54 ;
     RECT  98.595 160.43 98.755 160.54 ;
     RECT  118.855 160.42 118.965 160.54 ;
     RECT  1.985 160.395 2.155 160.565 ;
     RECT  2.72 160.395 2.89 160.565 ;
     RECT  6.585 160.395 6.755 160.565 ;
     RECT  11.46 160.395 11.63 160.565 ;
     RECT  15.785 160.395 15.955 160.565 ;
     RECT  16.245 160.395 16.415 160.565 ;
     RECT  23.145 160.395 23.315 160.565 ;
     RECT  30.505 160.395 30.675 160.565 ;
     RECT  35.565 160.395 35.735 160.565 ;
     RECT  37.86 160.395 38.03 160.565 ;
     RECT  40.625 160.395 40.795 160.565 ;
     RECT  43.66 160.395 43.83 160.565 ;
     RECT  47.525 160.395 47.695 160.565 ;
     RECT  51.67 160.395 51.84 160.565 ;
     RECT  55.16 160.395 55.33 160.565 ;
     RECT  57.46 160.395 57.63 160.565 ;
     RECT  61.325 160.395 61.495 160.565 ;
     RECT  62.52 160.395 62.69 160.565 ;
     RECT  68.96 160.395 69.13 160.565 ;
     RECT  70.985 160.395 71.155 160.565 ;
     RECT  73.1 160.395 73.27 160.565 ;
     RECT  76.965 160.395 77.135 160.565 ;
     RECT  78.62 160.395 78.79 160.565 ;
     RECT  82.945 160.395 83.115 160.565 ;
     RECT  85.06 160.395 85.23 160.565 ;
     RECT  88.925 160.395 89.095 160.565 ;
     RECT  90.765 160.395 90.935 160.565 ;
     RECT  92.88 160.395 93.05 160.565 ;
     RECT  98.125 160.395 98.295 160.565 ;
     RECT  100.24 160.395 100.41 160.565 ;
     RECT  104.105 160.395 104.275 160.565 ;
     RECT  106.68 160.395 106.85 160.565 ;
     RECT  111.465 160.535 111.635 160.565 ;
     RECT  113.305 160.395 113.475 160.565 ;
     RECT  47.97 160.43 48.19 160.6 ;
     RECT  15.325 160.8 15.495 161.325 ;
     RECT  42.925 160.8 43.095 161.325 ;
     RECT  70.525 160.8 70.695 161.325 ;
     RECT  98.125 160.8 98.295 161.325 ;
     RECT  29.125 165.075 29.295 165.6 ;
     RECT  56.725 165.075 56.895 165.6 ;
     RECT  84.325 165.075 84.495 165.6 ;
     RECT  111.925 165.075 112.095 165.6 ;
     RECT  1.535 165.86 1.695 165.865 ;
     RECT  1.52 165.865 1.695 165.97 ;
     RECT  7.055 165.86 7.215 165.97 ;
     RECT  15.335 165.86 15.495 165.97 ;
     RECT  28.215 165.86 28.375 165.97 ;
     RECT  55.815 165.86 55.975 165.97 ;
     RECT  57.195 165.86 57.355 165.97 ;
     RECT  63.635 165.86 63.795 165.97 ;
     RECT  70.97 165.8 71.19 165.97 ;
     RECT  96.295 165.86 96.455 165.97 ;
     RECT  119.755 165.86 119.915 165.97 ;
     RECT  1.52 165.97 1.64 165.975 ;
     RECT  2.44 165.865 2.56 165.975 ;
     RECT  16.24 165.865 16.36 165.975 ;
     RECT  22.68 165.865 22.8 165.975 ;
     RECT  42.46 165.865 42.58 165.975 ;
     RECT  52.58 165.865 52.7 165.975 ;
     RECT  58.1 165.865 58.22 165.975 ;
     RECT  70.06 165.865 70.18 165.975 ;
     RECT  71.9 165.865 72.02 165.975 ;
     RECT  75.58 165.865 75.7 165.975 ;
     RECT  83.86 165.865 83.98 165.975 ;
     RECT  97.2 165.865 97.32 165.975 ;
     RECT  99.5 165.865 99.62 165.975 ;
     RECT  105.94 165.865 106.06 165.975 ;
     RECT  120.66 165.865 120.78 165.975 ;
     RECT  9.355 165.87 9.515 165.98 ;
     RECT  14.415 165.87 14.575 165.98 ;
     RECT  15.815 165.86 15.925 165.98 ;
     RECT  21.775 165.87 21.935 165.98 ;
     RECT  51.675 165.87 51.835 165.98 ;
     RECT  53.995 165.86 54.105 165.98 ;
     RECT  74.675 165.87 74.835 165.98 ;
     RECT  98.595 165.87 98.755 165.98 ;
     RECT  101.835 165.86 101.945 165.98 ;
     RECT  118.855 165.86 118.965 165.98 ;
     RECT  1.985 165.835 2.155 166.005 ;
     RECT  3.18 165.835 3.35 166.005 ;
     RECT  7.965 165.835 8.135 166.005 ;
     RECT  10.54 165.835 10.71 166.005 ;
     RECT  16.98 165.835 17.15 166.005 ;
     RECT  17.9 165.835 18.07 166.005 ;
     RECT  20.85 165.835 21.02 166.005 ;
     RECT  23.145 165.835 23.315 166.005 ;
     RECT  29.585 165.835 29.755 166.005 ;
     RECT  30.505 165.835 30.675 166.005 ;
     RECT  36.945 165.835 37.115 166.005 ;
     RECT  37.87 165.835 38.04 166.005 ;
     RECT  43.66 165.835 43.83 166.005 ;
     RECT  44.305 165.835 44.475 166.005 ;
     RECT  47.8 165.835 47.97 166.005 ;
     RECT  53.045 165.835 53.215 166.005 ;
     RECT  58.57 165.835 58.74 166.005 ;
     RECT  60.405 165.835 60.575 166.005 ;
     RECT  64.545 165.835 64.715 166.005 ;
     RECT  72.365 165.835 72.535 166.005 ;
     RECT  76.045 165.835 76.215 166.005 ;
     RECT  80 165.835 80.17 166.005 ;
     RECT  83.405 165.835 83.575 166.005 ;
     RECT  84.785 165.835 84.955 166.005 ;
     RECT  87.085 165.835 87.255 166.005 ;
     RECT  90.765 165.835 90.935 166.005 ;
     RECT  92.42 165.835 92.59 166.005 ;
     RECT  94.445 165.835 94.615 166.005 ;
     RECT  97.94 165.835 98.11 166.005 ;
     RECT  100.24 165.835 100.41 166.005 ;
     RECT  103.65 165.835 103.82 166.005 ;
     RECT  104.11 165.835 104.28 166.005 ;
     RECT  106.68 165.835 106.85 166.005 ;
     RECT  108.245 165.835 108.415 166.005 ;
     RECT  110.82 165.835 110.99 166.005 ;
     RECT  112.385 165.835 112.555 166.005 ;
     RECT  114.96 165.835 115.13 166.005 ;
     RECT  15.325 166.24 15.495 166.765 ;
     RECT  42.925 166.24 43.095 166.765 ;
     RECT  70.525 166.24 70.695 166.765 ;
     RECT  98.125 166.24 98.295 166.765 ;
     RECT  29.125 170.515 29.295 171.04 ;
     RECT  56.725 170.515 56.895 171.04 ;
     RECT  84.325 170.515 84.495 171.04 ;
     RECT  111.925 170.515 112.095 171.04 ;
     RECT  1.535 171.3 1.695 171.305 ;
     RECT  1.52 171.305 1.695 171.41 ;
     RECT  23.615 171.3 23.775 171.41 ;
     RECT  59.035 171.3 59.195 171.41 ;
     RECT  112.395 171.3 112.555 171.41 ;
     RECT  1.52 171.41 1.64 171.415 ;
     RECT  2.44 171.305 2.56 171.415 ;
     RECT  24.52 171.305 24.64 171.415 ;
     RECT  44.3 171.305 44.42 171.415 ;
     RECT  70.98 171.305 71.1 171.415 ;
     RECT  78.8 171.305 78.92 171.415 ;
     RECT  83.86 171.305 83.98 171.415 ;
     RECT  84.78 171.305 84.9 171.415 ;
     RECT  120.66 171.305 120.78 171.415 ;
     RECT  9.375 171.3 9.485 171.42 ;
     RECT  15.795 171.31 15.955 171.42 ;
     RECT  21.795 171.3 21.905 171.42 ;
     RECT  29.615 171.3 29.725 171.42 ;
     RECT  41.115 171.3 41.225 171.42 ;
     RECT  43.395 171.31 43.555 171.42 ;
     RECT  50.775 171.3 50.885 171.42 ;
     RECT  57.215 171.3 57.325 171.42 ;
     RECT  59.515 171.3 59.625 171.42 ;
     RECT  68.715 171.3 68.825 171.42 ;
     RECT  1.985 171.275 2.155 171.445 ;
     RECT  3.18 171.275 3.35 171.445 ;
     RECT  7.045 171.275 7.215 171.445 ;
     RECT  11.46 171.275 11.63 171.445 ;
     RECT  14.405 171.275 14.575 171.445 ;
     RECT  16.705 171.275 16.875 171.445 ;
     RECT  24.065 171.275 24.235 171.445 ;
     RECT  25.26 171.275 25.43 171.445 ;
     RECT  31.425 171.275 31.595 171.445 ;
     RECT  38.79 171.275 38.96 171.445 ;
     RECT  44.765 171.275 44.935 171.445 ;
     RECT  46.15 171.275 46.32 171.445 ;
     RECT  52.125 171.275 52.295 171.445 ;
     RECT  52.86 171.275 53.03 171.445 ;
     RECT  60.22 171.275 60.39 171.445 ;
     RECT  61.325 171.275 61.495 171.445 ;
     RECT  64.085 171.275 64.255 171.445 ;
     RECT  71.445 171.275 71.615 171.445 ;
     RECT  71.72 171.275 71.89 171.445 ;
     RECT  75.86 171.275 76.03 171.445 ;
     RECT  79.265 171.275 79.435 171.445 ;
     RECT  79.73 171.275 79.9 171.445 ;
     RECT  85.245 171.275 85.415 171.445 ;
     RECT  86.63 171.275 86.8 171.445 ;
     RECT  90.765 171.275 90.935 171.445 ;
     RECT  92.61 171.275 92.78 171.445 ;
     RECT  96.75 171.275 96.92 171.445 ;
     RECT  98.585 171.275 98.755 171.445 ;
     RECT  100.885 171.275 101.055 171.445 ;
     RECT  104.565 171.275 104.735 171.445 ;
     RECT  106.22 171.275 106.39 171.445 ;
     RECT  110.085 171.275 110.255 171.445 ;
     RECT  113.305 171.275 113.475 171.445 ;
     RECT  113.765 171.275 113.935 171.445 ;
     RECT  15.325 171.68 15.495 172.205 ;
     RECT  42.925 171.68 43.095 172.205 ;
     RECT  70.525 171.68 70.695 172.205 ;
     RECT  98.125 171.68 98.295 172.205 ;
     RECT  29.125 175.955 29.295 176.48 ;
     RECT  56.725 175.955 56.895 176.48 ;
     RECT  84.325 175.955 84.495 176.48 ;
     RECT  111.925 175.955 112.095 176.48 ;
     RECT  1.535 176.74 1.695 176.745 ;
     RECT  66.395 176.74 66.555 176.745 ;
     RECT  1.52 176.745 1.695 176.85 ;
     RECT  6.595 176.74 6.755 176.85 ;
     RECT  42.935 176.74 43.095 176.85 ;
     RECT  55.815 176.74 55.975 176.85 ;
     RECT  66.38 176.745 66.555 176.85 ;
     RECT  111.015 176.74 111.175 176.85 ;
     RECT  1.52 176.85 1.64 176.855 ;
     RECT  24.06 176.745 24.18 176.855 ;
     RECT  24.52 176.745 24.64 176.855 ;
     RECT  43.84 176.745 43.96 176.855 ;
     RECT  50.28 176.745 50.4 176.855 ;
     RECT  66.38 176.85 66.5 176.855 ;
     RECT  67.3 176.745 67.42 176.855 ;
     RECT  120.66 176.745 120.78 176.855 ;
     RECT  9.375 176.74 9.485 176.86 ;
     RECT  15.795 176.75 15.955 176.86 ;
     RECT  29.615 176.74 29.725 176.86 ;
     RECT  40.195 176.74 40.305 176.86 ;
     RECT  42.015 176.75 42.175 176.86 ;
     RECT  43.415 176.74 43.525 176.86 ;
     RECT  45.235 176.75 45.395 176.86 ;
     RECT  64.575 176.74 64.685 176.86 ;
     RECT  76.975 176.75 77.135 176.86 ;
     RECT  118.855 176.74 118.965 176.86 ;
     RECT  1.985 176.715 2.155 176.885 ;
     RECT  2.72 176.715 2.89 176.885 ;
     RECT  7.505 176.715 7.675 176.885 ;
     RECT  11.46 176.715 11.63 176.885 ;
     RECT  16.705 176.715 16.875 176.885 ;
     RECT  17.165 176.715 17.335 176.885 ;
     RECT  24.8 176.715 24.97 176.885 ;
     RECT  25.26 176.715 25.43 176.885 ;
     RECT  28.67 176.715 28.84 176.885 ;
     RECT  31.425 176.715 31.595 176.885 ;
     RECT  32.805 176.715 32.975 176.885 ;
     RECT  39.06 176.715 39.23 176.885 ;
     RECT  44.305 176.715 44.475 176.885 ;
     RECT  46.42 176.715 46.59 176.885 ;
     RECT  50.745 176.715 50.915 176.885 ;
     RECT  51.94 176.715 52.11 176.885 ;
     RECT  57.185 176.715 57.355 176.885 ;
     RECT  60.68 176.715 60.85 176.885 ;
     RECT  66.845 176.715 67.015 176.885 ;
     RECT  67.765 176.715 67.935 176.885 ;
     RECT  71.26 176.715 71.43 176.885 ;
     RECT  75.125 176.715 75.295 176.885 ;
     RECT  77.885 176.715 78.055 176.885 ;
     RECT  84.785 176.715 84.955 176.885 ;
     RECT  87.085 176.715 87.255 176.885 ;
     RECT  92.145 176.715 92.315 176.885 ;
     RECT  94.445 176.715 94.615 176.885 ;
     RECT  98.86 176.715 99.03 176.885 ;
     RECT  99.505 176.715 99.675 176.885 ;
     RECT  102.73 176.715 102.9 176.885 ;
     RECT  105.485 176.715 105.655 176.885 ;
     RECT  107.14 176.715 107.31 176.885 ;
     RECT  112.39 176.715 112.56 176.885 ;
     RECT  114.96 176.715 115.13 176.885 ;
     RECT  117.26 176.715 117.43 176.885 ;
     RECT  15.325 177.12 15.495 177.645 ;
     RECT  42.925 177.12 43.095 177.645 ;
     RECT  70.525 177.12 70.695 177.645 ;
     RECT  98.125 177.12 98.295 177.645 ;
     RECT  29.125 181.395 29.295 181.92 ;
     RECT  56.725 181.395 56.895 181.92 ;
     RECT  84.325 181.395 84.495 181.92 ;
     RECT  111.925 181.395 112.095 181.92 ;
     RECT  1.535 182.18 1.695 182.185 ;
     RECT  16.705 182.155 16.875 182.185 ;
     RECT  1.52 182.185 1.695 182.29 ;
     RECT  8.435 182.18 8.595 182.29 ;
     RECT  27.755 182.18 27.915 182.29 ;
     RECT  29.595 182.18 29.755 182.29 ;
     RECT  55.355 182.18 55.515 182.29 ;
     RECT  93.075 182.18 93.235 182.29 ;
     RECT  102.275 182.18 102.435 182.29 ;
     RECT  111.015 182.18 111.175 182.29 ;
     RECT  1.52 182.29 1.64 182.295 ;
     RECT  16.7 182.185 16.875 182.295 ;
     RECT  28.66 182.185 28.78 182.295 ;
     RECT  56.26 182.185 56.38 182.295 ;
     RECT  68.68 182.185 68.8 182.295 ;
     RECT  83.4 182.185 83.52 182.295 ;
     RECT  87.54 182.185 87.66 182.295 ;
     RECT  97.66 182.185 97.78 182.295 ;
     RECT  103.18 182.185 103.3 182.295 ;
     RECT  112.84 182.185 112.96 182.295 ;
     RECT  120.66 182.185 120.78 182.295 ;
     RECT  6.615 182.18 6.725 182.3 ;
     RECT  15.795 182.19 15.955 182.3 ;
     RECT  25.935 182.18 26.045 182.3 ;
     RECT  69.615 182.19 69.775 182.3 ;
     RECT  75.135 182.19 75.295 182.3 ;
     RECT  95.855 182.18 95.965 182.3 ;
     RECT  102.755 182.18 102.865 182.3 ;
     RECT  104.575 182.19 104.735 182.3 ;
     RECT  1.985 182.155 2.155 182.325 ;
     RECT  2.72 182.155 2.89 182.325 ;
     RECT  9.345 182.155 9.515 182.325 ;
     RECT  11.46 182.155 11.63 182.325 ;
     RECT  16.705 182.295 16.875 182.325 ;
     RECT  17.44 182.155 17.61 182.325 ;
     RECT  21.305 182.155 21.475 182.325 ;
     RECT  30.78 182.155 30.95 182.325 ;
     RECT  30.965 182.155 31.135 182.325 ;
     RECT  34.645 182.155 34.815 182.325 ;
     RECT  38.33 182.155 38.5 182.325 ;
     RECT  43.385 182.155 43.555 182.325 ;
     RECT  43.845 182.155 44.015 182.325 ;
     RECT  51.48 182.155 51.65 182.325 ;
     RECT  53.045 182.155 53.215 182.325 ;
     RECT  57.46 182.155 57.63 182.325 ;
     RECT  61.325 182.155 61.495 182.325 ;
     RECT  62.245 182.155 62.415 182.325 ;
     RECT  69.42 182.155 69.59 182.325 ;
     RECT  71.26 182.155 71.43 182.325 ;
     RECT  73.285 182.155 73.455 182.325 ;
     RECT  76.045 182.155 76.215 182.325 ;
     RECT  80.645 182.155 80.815 182.325 ;
     RECT  83.865 182.155 84.035 182.325 ;
     RECT  85.06 182.155 85.23 182.325 ;
     RECT  88.28 182.155 88.45 182.325 ;
     RECT  89.2 182.155 89.37 182.325 ;
     RECT  92.145 182.155 92.315 182.325 ;
     RECT  93.99 182.155 94.16 182.325 ;
     RECT  98.13 182.155 98.3 182.325 ;
     RECT  98.86 182.155 99.03 182.325 ;
     RECT  103.645 182.155 103.815 182.325 ;
     RECT  105.485 182.155 105.655 182.325 ;
     RECT  112.66 182.155 112.83 182.325 ;
     RECT  113.305 182.155 113.475 182.325 ;
     RECT  116.8 182.155 116.97 182.325 ;
     RECT  15.325 182.56 15.495 183.085 ;
     RECT  42.925 182.56 43.095 183.085 ;
     RECT  70.525 182.56 70.695 183.085 ;
     RECT  98.125 182.56 98.295 183.085 ;
     RECT  29.125 186.835 29.295 187.36 ;
     RECT  56.725 186.835 56.895 187.36 ;
     RECT  84.325 186.835 84.495 187.36 ;
     RECT  111.925 186.835 112.095 187.36 ;
     RECT  55.355 187.62 55.515 187.625 ;
     RECT  3.375 187.62 3.535 187.73 ;
     RECT  36.495 187.62 36.655 187.73 ;
     RECT  50.295 187.62 50.455 187.73 ;
     RECT  55.34 187.625 55.515 187.73 ;
     RECT  4.28 187.625 4.4 187.735 ;
     RECT  21.3 187.625 21.42 187.735 ;
     RECT  37.4 187.625 37.52 187.735 ;
     RECT  50.74 187.625 50.86 187.735 ;
     RECT  55.34 187.73 55.46 187.735 ;
     RECT  56.26 187.625 56.38 187.735 ;
     RECT  70.06 187.625 70.18 187.735 ;
     RECT  71.9 187.625 72.02 187.735 ;
     RECT  77.88 187.625 78 187.735 ;
     RECT  91.68 187.625 91.8 187.735 ;
     RECT  97.66 187.625 97.78 187.735 ;
     RECT  111.46 187.625 111.58 187.735 ;
     RECT  120.66 187.625 120.78 187.735 ;
     RECT  1.555 187.62 1.665 187.74 ;
     RECT  19.495 187.62 19.605 187.74 ;
     RECT  27.295 187.63 27.455 187.74 ;
     RECT  34.675 187.62 34.785 187.74 ;
     RECT  68.255 187.62 68.365 187.74 ;
     RECT  70.995 187.63 71.155 187.74 ;
     RECT  82.515 187.62 82.625 187.74 ;
     RECT  84.815 187.62 84.925 187.74 ;
     RECT  90.775 187.63 90.935 187.74 ;
     RECT  95.855 187.62 95.965 187.74 ;
     RECT  1.8 187.595 1.97 187.765 ;
     RECT  4.745 187.595 4.915 187.765 ;
     RECT  5.665 187.595 5.835 187.765 ;
     RECT  12.105 187.595 12.275 187.765 ;
     RECT  15.785 187.595 15.955 187.765 ;
     RECT  21.765 187.595 21.935 187.765 ;
     RECT  23.42 187.595 23.59 187.765 ;
     RECT  28.205 187.595 28.375 187.765 ;
     RECT  29.59 187.595 29.76 187.765 ;
     RECT  35.565 187.595 35.735 187.765 ;
     RECT  37.87 187.595 38.04 187.765 ;
     RECT  42.925 187.595 43.095 187.765 ;
     RECT  43.385 187.595 43.555 187.765 ;
     RECT  51.48 187.595 51.65 187.765 ;
     RECT  55.81 187.595 55.98 187.765 ;
     RECT  57.19 187.595 57.36 187.765 ;
     RECT  60.865 187.595 61.035 187.765 ;
     RECT  64.36 187.595 64.53 187.765 ;
     RECT  70.525 187.595 70.695 187.765 ;
     RECT  72.365 187.595 72.535 187.765 ;
     RECT  78.62 187.595 78.79 187.765 ;
     RECT  79.725 187.595 79.895 187.765 ;
     RECT  86.625 187.595 86.795 187.765 ;
     RECT  87.09 187.595 87.26 187.765 ;
     RECT  92.15 187.595 92.32 187.765 ;
     RECT  93.99 187.595 94.16 187.765 ;
     RECT  96.745 187.595 96.915 187.765 ;
     RECT  98.585 187.595 98.755 187.765 ;
     RECT  102.265 187.595 102.435 187.765 ;
     RECT  104.105 187.595 104.275 187.765 ;
     RECT  109.9 187.595 110.07 187.765 ;
     RECT  112.66 187.595 112.83 187.765 ;
     RECT  113.765 187.595 113.935 187.765 ;
     RECT  116.8 187.595 116.97 187.765 ;
     RECT  15.325 188 15.495 188.525 ;
     RECT  42.925 188 43.095 188.525 ;
     RECT  70.525 188 70.695 188.525 ;
     RECT  98.125 188 98.295 188.525 ;
     RECT  29.125 192.275 29.295 192.8 ;
     RECT  56.725 192.275 56.895 192.8 ;
     RECT  84.325 192.275 84.495 192.8 ;
     RECT  111.925 192.275 112.095 192.8 ;
     RECT  32.345 193.035 32.515 193.065 ;
     RECT  1.52 193.065 1.64 193.07 ;
     RECT  31.435 193.06 31.595 193.17 ;
     RECT  48.455 193.06 48.615 193.17 ;
     RECT  64.095 193.06 64.255 193.17 ;
     RECT  88.935 193.06 89.095 193.17 ;
     RECT  97.675 193.06 97.835 193.17 ;
     RECT  120.215 193.06 120.375 193.17 ;
     RECT  1.52 193.07 1.695 193.175 ;
     RECT  2.44 193.065 2.56 193.175 ;
     RECT  32.34 193.065 32.515 193.175 ;
     RECT  42.46 193.065 42.58 193.175 ;
     RECT  44.3 193.065 44.42 193.175 ;
     RECT  65 193.065 65.12 193.175 ;
     RECT  89.84 193.065 89.96 193.175 ;
     RECT  1.535 193.175 1.695 193.18 ;
     RECT  7.055 193.07 7.215 193.18 ;
     RECT  9.375 193.06 9.485 193.18 ;
     RECT  15.355 193.06 15.465 193.18 ;
     RECT  24.075 193.07 24.235 193.18 ;
     RECT  29.615 193.06 29.725 193.18 ;
     RECT  39.735 193.06 39.845 193.18 ;
     RECT  41.555 193.07 41.715 193.18 ;
     RECT  43.395 193.07 43.555 193.18 ;
     RECT  46.635 193.06 46.745 193.18 ;
     RECT  48.935 193.06 49.045 193.18 ;
     RECT  62.275 193.06 62.385 193.18 ;
     RECT  67.795 193.06 67.905 193.18 ;
     RECT  91.255 193.06 91.365 193.18 ;
     RECT  93.075 193.07 93.235 193.18 ;
     RECT  1.985 193.035 2.155 193.205 ;
     RECT  3.18 193.035 3.35 193.205 ;
     RECT  7.965 193.035 8.135 193.205 ;
     RECT  11.19 193.035 11.36 193.205 ;
     RECT  16.06 193.035 16.23 193.205 ;
     RECT  17.44 193.035 17.61 193.205 ;
     RECT  20.2 193.035 20.37 193.205 ;
     RECT  21.305 193.035 21.475 193.205 ;
     RECT  24.985 193.035 25.155 193.205 ;
     RECT  25.26 193.035 25.43 193.205 ;
     RECT  32.345 193.175 32.515 193.205 ;
     RECT  32.805 193.035 32.975 193.205 ;
     RECT  42.74 193.035 42.91 193.205 ;
     RECT  45.04 193.035 45.21 193.205 ;
     RECT  49.365 193.035 49.535 193.205 ;
     RECT  50.745 193.035 50.915 193.205 ;
     RECT  57.19 193.035 57.36 193.205 ;
     RECT  60.405 193.035 60.575 193.205 ;
     RECT  65.74 193.035 65.91 193.205 ;
     RECT  69.605 193.035 69.775 193.205 ;
     RECT  71.26 193.035 71.43 193.205 ;
     RECT  75.4 193.035 75.57 193.205 ;
     RECT  76.965 193.035 77.135 193.205 ;
     RECT  79.54 193.035 79.71 193.205 ;
     RECT  83.68 193.035 83.85 193.205 ;
     RECT  85.06 193.035 85.23 193.205 ;
     RECT  87.545 193.035 87.715 193.205 ;
     RECT  90.305 193.035 90.475 193.205 ;
     RECT  94.26 193.035 94.43 193.205 ;
     RECT  98.59 193.035 98.76 193.205 ;
     RECT  102.265 193.035 102.435 193.205 ;
     RECT  103.46 193.035 103.63 193.205 ;
     RECT  107.33 193.035 107.5 193.205 ;
     RECT  109.9 193.035 110.07 193.205 ;
     RECT  112.385 193.035 112.555 193.205 ;
     RECT  114.04 193.035 114.21 193.205 ;
     RECT  116.34 193.035 116.51 193.205 ;
     RECT  117.905 193.035 118.075 193.205 ;
     RECT  15.325 193.44 15.495 193.965 ;
     RECT  42.925 193.44 43.095 193.965 ;
     RECT  70.525 193.44 70.695 193.965 ;
     RECT  98.125 193.44 98.295 193.965 ;
     RECT  29.125 197.715 29.295 198.24 ;
     RECT  56.725 197.715 56.895 198.24 ;
     RECT  84.325 197.715 84.495 198.24 ;
     RECT  111.925 197.715 112.095 198.24 ;
     RECT  1.555 198.5 1.665 198.505 ;
     RECT  28.215 198.5 28.375 198.61 ;
     RECT  61.335 198.5 61.495 198.61 ;
     RECT  71.455 198.5 71.615 198.61 ;
     RECT  91.695 198.5 91.855 198.61 ;
     RECT  103.655 198.5 103.815 198.61 ;
     RECT  119.755 198.5 119.915 198.61 ;
     RECT  1.52 198.505 1.665 198.615 ;
     RECT  11.18 198.505 11.3 198.615 ;
     RECT  14.86 198.505 14.98 198.615 ;
     RECT  70.06 198.505 70.18 198.615 ;
     RECT  83.86 198.505 83.98 198.615 ;
     RECT  84.78 198.505 84.9 198.615 ;
     RECT  120.66 198.505 120.78 198.615 ;
     RECT  1.555 198.615 1.665 198.62 ;
     RECT  9.375 198.5 9.485 198.62 ;
     RECT  19.935 198.51 20.095 198.62 ;
     RECT  26.395 198.5 26.505 198.62 ;
     RECT  37.875 198.51 38.035 198.62 ;
     RECT  47.535 198.51 47.695 198.62 ;
     RECT  68.255 198.5 68.365 198.62 ;
     RECT  69.635 198.5 69.745 198.62 ;
     RECT  76.535 198.5 76.645 198.62 ;
     RECT  89.875 198.5 89.985 198.62 ;
     RECT  1.985 198.475 2.155 198.645 ;
     RECT  3.64 198.475 3.81 198.645 ;
     RECT  7.505 198.475 7.675 198.645 ;
     RECT  11.645 198.475 11.815 198.645 ;
     RECT  16.06 198.475 16.23 198.645 ;
     RECT  19.005 198.475 19.175 198.645 ;
     RECT  20.845 198.475 21.015 198.645 ;
     RECT  29.86 198.475 30.03 198.645 ;
     RECT  30.505 198.475 30.675 198.645 ;
     RECT  34 198.475 34.17 198.645 ;
     RECT  38.14 198.475 38.31 198.645 ;
     RECT  39.06 198.475 39.23 198.645 ;
     RECT  42.005 198.475 42.175 198.645 ;
     RECT  43.66 198.475 43.83 198.645 ;
     RECT  48.72 198.475 48.89 198.645 ;
     RECT  49.365 198.475 49.535 198.645 ;
     RECT  52.86 198.475 53.03 198.645 ;
     RECT  57 198.475 57.17 198.645 ;
     RECT  57.46 198.475 57.63 198.645 ;
     RECT  60.865 198.475 61.035 198.645 ;
     RECT  62.245 198.475 62.415 198.645 ;
     RECT  70.985 198.475 71.155 198.645 ;
     RECT  72.64 198.475 72.81 198.645 ;
     RECT  78.345 198.475 78.515 198.645 ;
     RECT  82.03 198.475 82.2 198.645 ;
     RECT  85.25 198.475 85.42 198.645 ;
     RECT  86.625 198.475 86.795 198.645 ;
     RECT  92.605 198.475 92.775 198.645 ;
     RECT  94.26 198.475 94.43 198.645 ;
     RECT  98.585 198.475 98.755 198.645 ;
     RECT  99.965 198.475 100.135 198.645 ;
     RECT  104.565 198.475 104.735 198.645 ;
     RECT  105.945 198.475 106.115 198.645 ;
     RECT  112.385 198.475 112.555 198.645 ;
     RECT  113.58 198.475 113.75 198.645 ;
     RECT  117.445 198.475 117.615 198.645 ;
     RECT  15.325 198.88 15.495 199.405 ;
     RECT  42.925 198.88 43.095 199.405 ;
     RECT  70.525 198.88 70.695 199.405 ;
     RECT  98.125 198.88 98.295 199.405 ;
     RECT  29.125 203.155 29.295 203.68 ;
     RECT  56.725 203.155 56.895 203.68 ;
     RECT  84.325 203.155 84.495 203.68 ;
     RECT  111.925 203.155 112.095 203.68 ;
     RECT  5.675 203.94 5.835 204.05 ;
     RECT  22.695 203.94 22.855 204.05 ;
     RECT  28.215 203.94 28.375 204.05 ;
     RECT  29.595 203.94 29.755 204.05 ;
     RECT  45.695 203.94 45.855 204.05 ;
     RECT  55.815 203.94 55.975 204.05 ;
     RECT  71.455 203.94 71.615 204.05 ;
     RECT  106.415 203.94 106.575 204.05 ;
     RECT  2.44 203.945 2.56 204.055 ;
     RECT  6.58 203.945 6.7 204.055 ;
     RECT  23.6 203.945 23.72 204.055 ;
     RECT  30.5 203.945 30.62 204.055 ;
     RECT  43.38 203.945 43.5 204.055 ;
     RECT  71.9 203.945 72.02 204.055 ;
     RECT  83.86 203.945 83.98 204.055 ;
     RECT  104.56 203.945 104.68 204.055 ;
     RECT  111.46 203.945 111.58 204.055 ;
     RECT  113.3 203.945 113.42 204.055 ;
     RECT  120.66 203.945 120.78 204.055 ;
     RECT  1.535 203.95 1.695 204.06 ;
     RECT  14.415 203.95 14.575 204.06 ;
     RECT  20.875 203.94 20.985 204.06 ;
     RECT  53.995 203.94 54.105 204.06 ;
     RECT  69.635 203.94 69.745 204.06 ;
     RECT  70.995 203.95 71.155 204.06 ;
     RECT  93.095 203.94 93.205 204.06 ;
     RECT  103.655 203.95 103.815 204.06 ;
     RECT  117.935 203.94 118.045 204.06 ;
     RECT  119.755 203.95 119.915 204.06 ;
     RECT  1.8 203.915 1.97 204.085 ;
     RECT  2.905 203.915 3.075 204.085 ;
     RECT  7.045 203.915 7.215 204.085 ;
     RECT  10.54 203.915 10.71 204.085 ;
     RECT  15.785 203.915 15.955 204.085 ;
     RECT  16.98 203.915 17.15 204.085 ;
     RECT  23.42 203.915 23.59 204.085 ;
     RECT  24.34 203.915 24.51 204.085 ;
     RECT  27.56 203.915 27.73 204.085 ;
     RECT  30.965 203.915 31.135 204.085 ;
     RECT  31.7 203.915 31.87 204.085 ;
     RECT  35.565 203.915 35.735 204.085 ;
     RECT  38.325 203.915 38.495 204.085 ;
     RECT  43.845 203.915 44.015 204.085 ;
     RECT  46.605 203.915 46.775 204.085 ;
     RECT  53.505 203.915 53.675 204.085 ;
     RECT  57.19 203.915 57.36 204.085 ;
     RECT  63.165 203.915 63.335 204.085 ;
     RECT  65.74 203.915 65.91 204.085 ;
     RECT  72.365 203.915 72.535 204.085 ;
     RECT  79.725 203.915 79.895 204.085 ;
     RECT  80 203.915 80.17 204.085 ;
     RECT  85.06 203.915 85.23 204.085 ;
     RECT  87.085 203.915 87.255 204.085 ;
     RECT  89.2 203.915 89.37 204.085 ;
     RECT  94.445 203.915 94.615 204.085 ;
     RECT  94.905 203.915 95.075 204.085 ;
     RECT  98.59 203.915 98.76 204.085 ;
     RECT  102.54 203.915 102.71 204.085 ;
     RECT  105.3 203.915 105.47 204.085 ;
     RECT  107.6 203.915 107.77 204.085 ;
     RECT  109.44 203.915 109.61 204.085 ;
     RECT  112.39 203.915 112.56 204.085 ;
     RECT  114.04 203.915 114.21 204.085 ;
     RECT  117.26 203.915 117.43 204.085 ;
     RECT  15.325 204.32 15.495 204.845 ;
     RECT  42.925 204.32 43.095 204.845 ;
     RECT  70.525 204.32 70.695 204.845 ;
     RECT  98.125 204.32 98.295 204.845 ;
     RECT  29.125 208.595 29.295 209.12 ;
     RECT  56.725 208.595 56.895 209.12 ;
     RECT  84.325 208.595 84.495 209.12 ;
     RECT  111.925 208.595 112.095 209.12 ;
     RECT  1.555 209.38 1.665 209.385 ;
     RECT  33.735 209.38 33.895 209.49 ;
     RECT  55.815 209.38 55.975 209.49 ;
     RECT  66.855 209.38 67.015 209.49 ;
     RECT  78.815 209.38 78.975 209.49 ;
     RECT  97.675 209.38 97.835 209.49 ;
     RECT  111.015 209.38 111.175 209.49 ;
     RECT  120.215 209.38 120.375 209.49 ;
     RECT  1.52 209.385 1.665 209.495 ;
     RECT  17.62 209.385 17.74 209.495 ;
     RECT  28.66 209.385 28.78 209.495 ;
     RECT  34.64 209.385 34.76 209.495 ;
     RECT  37.86 209.385 37.98 209.495 ;
     RECT  45.22 209.385 45.34 209.495 ;
     RECT  59.02 209.385 59.14 209.495 ;
     RECT  79.72 209.385 79.84 209.495 ;
     RECT  84.32 209.385 84.44 209.495 ;
     RECT  92.14 209.385 92.26 209.495 ;
     RECT  111.46 209.385 111.58 209.495 ;
     RECT  112.38 209.385 112.5 209.495 ;
     RECT  1.555 209.495 1.665 209.5 ;
     RECT  3.375 209.39 3.535 209.5 ;
     RECT  13.515 209.38 13.625 209.5 ;
     RECT  15.815 209.38 15.925 209.5 ;
     RECT  26.855 209.38 26.965 209.5 ;
     RECT  29.595 209.39 29.755 209.5 ;
     RECT  43.415 209.38 43.525 209.5 ;
     RECT  57.215 209.38 57.325 209.5 ;
     RECT  69.615 209.39 69.775 209.5 ;
     RECT  76.995 209.38 77.105 209.5 ;
     RECT  83.415 209.39 83.575 209.5 ;
     RECT  89.855 209.39 90.015 209.5 ;
     RECT  109.655 209.38 109.765 209.5 ;
     RECT  1.985 209.355 2.155 209.525 ;
     RECT  4.285 209.355 4.455 209.525 ;
     RECT  9.62 209.355 9.79 209.525 ;
     RECT  15.325 209.355 15.495 209.525 ;
     RECT  18.36 209.355 18.53 209.525 ;
     RECT  22.225 209.355 22.395 209.525 ;
     RECT  22.96 209.355 23.13 209.525 ;
     RECT  29.86 209.355 30.03 209.525 ;
     RECT  30.505 209.355 30.675 209.525 ;
     RECT  35.105 209.355 35.275 209.525 ;
     RECT  38.33 209.355 38.5 209.525 ;
     RECT  44.305 209.355 44.475 209.525 ;
     RECT  45.96 209.355 46.13 209.525 ;
     RECT  50.1 209.355 50.27 209.525 ;
     RECT  51.94 209.355 52.11 209.525 ;
     RECT  53.965 209.355 54.135 209.525 ;
     RECT  59.485 209.355 59.655 209.525 ;
     RECT  61.6 209.355 61.77 209.525 ;
     RECT  65.74 209.355 65.91 209.525 ;
     RECT  67.765 209.355 67.935 209.525 ;
     RECT  71.26 209.355 71.43 209.525 ;
     RECT  75.4 209.355 75.57 209.525 ;
     RECT  79.54 209.355 79.71 209.525 ;
     RECT  80.46 209.355 80.63 209.525 ;
     RECT  84.79 209.355 84.96 209.525 ;
     RECT  89.39 209.355 89.56 209.525 ;
     RECT  90.765 209.355 90.935 209.525 ;
     RECT  92.61 209.355 92.78 209.525 ;
     RECT  98.59 209.355 98.76 209.525 ;
     RECT  98.86 209.355 99.03 209.525 ;
     RECT  101.345 209.355 101.515 209.525 ;
     RECT  102.265 209.355 102.435 209.525 ;
     RECT  103 209.355 103.17 209.525 ;
     RECT  107.14 209.355 107.31 209.525 ;
     RECT  111.925 209.355 112.095 209.525 ;
     RECT  112.845 209.355 113.015 209.525 ;
     RECT  15.325 209.76 15.495 210.285 ;
     RECT  42.925 209.76 43.095 210.285 ;
     RECT  70.525 209.76 70.695 210.285 ;
     RECT  98.125 209.76 98.295 210.285 ;
     RECT  29.125 214.035 29.295 214.56 ;
     RECT  56.725 214.035 56.895 214.56 ;
     RECT  84.325 214.035 84.495 214.56 ;
     RECT  111.925 214.035 112.095 214.56 ;
     RECT  46.605 214.795 46.775 214.825 ;
     RECT  61.355 214.82 61.465 214.825 ;
     RECT  97.675 214.82 97.835 214.825 ;
     RECT  55.355 214.82 55.515 214.93 ;
     RECT  71.455 214.82 71.615 214.93 ;
     RECT  97.66 214.825 97.835 214.93 ;
     RECT  110.555 214.82 110.715 214.93 ;
     RECT  120.215 214.82 120.375 214.93 ;
     RECT  16.7 214.825 16.82 214.935 ;
     RECT  28.66 214.825 28.78 214.935 ;
     RECT  38.32 214.825 38.44 214.935 ;
     RECT  46.14 214.825 46.26 214.935 ;
     RECT  46.6 214.825 46.775 214.935 ;
     RECT  56.26 214.825 56.38 214.935 ;
     RECT  61.32 214.825 61.465 214.935 ;
     RECT  70.06 214.825 70.18 214.935 ;
     RECT  83.86 214.825 83.98 214.935 ;
     RECT  97.66 214.93 97.78 214.935 ;
     RECT  111.46 214.825 111.58 214.935 ;
     RECT  112.38 214.825 112.5 214.935 ;
     RECT  15.795 214.83 15.955 214.94 ;
     RECT  43.415 214.82 43.525 214.94 ;
     RECT  45.235 214.83 45.395 214.94 ;
     RECT  61.355 214.935 61.465 214.94 ;
     RECT  69.155 214.83 69.315 214.94 ;
     RECT  78.355 214.83 78.515 214.94 ;
     RECT  95.855 214.82 95.965 214.94 ;
     RECT  119.315 214.82 119.425 214.94 ;
     RECT  1.53 214.795 1.7 214.965 ;
     RECT  3.64 214.795 3.81 214.965 ;
     RECT  7.505 214.795 7.675 214.965 ;
     RECT  11.645 214.795 11.815 214.965 ;
     RECT  17.165 214.795 17.335 214.965 ;
     RECT  24.8 214.795 24.97 214.965 ;
     RECT  27.1 214.795 27.27 214.965 ;
     RECT  29.585 214.795 29.755 214.965 ;
     RECT  30.965 214.795 31.135 214.965 ;
     RECT  39.06 214.795 39.23 214.965 ;
     RECT  39.245 214.795 39.415 214.965 ;
     RECT  46.605 214.935 46.775 214.965 ;
     RECT  47.34 214.795 47.51 214.965 ;
     RECT  51.48 214.795 51.65 214.965 ;
     RECT  53.965 214.795 54.135 214.965 ;
     RECT  57.46 214.795 57.63 214.965 ;
     RECT  61.785 214.795 61.955 214.965 ;
     RECT  63.44 214.795 63.61 214.965 ;
     RECT  67.58 214.795 67.75 214.965 ;
     RECT  70.985 214.795 71.155 214.965 ;
     RECT  72.365 214.795 72.535 214.965 ;
     RECT  79.27 214.795 79.44 214.965 ;
     RECT  80 214.795 80.17 214.965 ;
     RECT  84.325 214.795 84.495 214.965 ;
     RECT  84.785 214.795 84.955 214.965 ;
     RECT  88.465 214.795 88.635 214.965 ;
     RECT  91.96 214.795 92.13 214.965 ;
     RECT  98.585 214.795 98.76 214.965 ;
     RECT  103.185 214.795 103.355 214.965 ;
     RECT  108.06 214.795 108.23 214.965 ;
     RECT  111.925 214.795 112.095 214.965 ;
     RECT  112.845 214.795 113.015 214.965 ;
     RECT  15.325 215.2 15.495 215.725 ;
     RECT  42.925 215.2 43.095 215.725 ;
     RECT  70.525 215.2 70.695 215.725 ;
     RECT  98.125 215.2 98.295 215.725 ;
     RECT  29.125 219.475 29.295 220 ;
     RECT  56.725 219.475 56.895 220 ;
     RECT  84.325 219.475 84.495 220 ;
     RECT  111.925 219.475 112.095 220 ;
     RECT  1.525 220.235 1.695 220.265 ;
     RECT  16.705 220.235 16.875 220.265 ;
     RECT  24.075 220.26 24.235 220.37 ;
     RECT  73.295 220.26 73.455 220.37 ;
     RECT  101.355 220.26 101.515 220.37 ;
     RECT  119.755 220.26 119.915 220.37 ;
     RECT  1.52 220.265 1.695 220.375 ;
     RECT  8.88 220.265 9 220.375 ;
     RECT  16.7 220.265 16.875 220.375 ;
     RECT  37.86 220.265 37.98 220.375 ;
     RECT  54.42 220.265 54.54 220.375 ;
     RECT  61.32 220.265 61.44 220.375 ;
     RECT  70.98 220.265 71.1 220.375 ;
     RECT  74.2 220.265 74.32 220.375 ;
     RECT  83.86 220.265 83.98 220.375 ;
     RECT  88.46 220.265 88.58 220.375 ;
     RECT  102.26 220.265 102.38 220.375 ;
     RECT  120.66 220.265 120.78 220.375 ;
     RECT  13.515 220.26 13.625 220.38 ;
     RECT  15.795 220.27 15.955 220.38 ;
     RECT  42.015 220.27 42.175 220.38 ;
     RECT  43.415 220.26 43.525 220.38 ;
     RECT  53.515 220.27 53.675 220.38 ;
     RECT  75.595 220.27 75.755 220.38 ;
     RECT  80.655 220.27 80.815 220.38 ;
     RECT  82.055 220.26 82.165 220.38 ;
     RECT  86.655 220.26 86.765 220.38 ;
     RECT  110.115 220.26 110.225 220.38 ;
     RECT  120.215 220.27 120.375 220.38 ;
     RECT  1.525 220.375 1.695 220.405 ;
     RECT  1.985 220.235 2.155 220.405 ;
     RECT  9.345 220.235 9.515 220.405 ;
     RECT  9.62 220.235 9.79 220.405 ;
     RECT  16.705 220.375 16.875 220.405 ;
     RECT  17.165 220.235 17.335 220.405 ;
     RECT  24.8 220.235 24.97 220.405 ;
     RECT  25.26 220.235 25.43 220.405 ;
     RECT  28.67 220.235 28.84 220.405 ;
     RECT  29.585 220.235 29.755 220.405 ;
     RECT  36.95 220.235 37.12 220.405 ;
     RECT  38.325 220.235 38.495 220.405 ;
     RECT  45.225 220.235 45.395 220.405 ;
     RECT  45.685 220.235 45.855 220.405 ;
     RECT  53.05 220.235 53.22 220.405 ;
     RECT  54.885 220.235 55.055 220.405 ;
     RECT  57.46 220.235 57.63 220.405 ;
     RECT  61.785 220.235 61.955 220.405 ;
     RECT  62.25 220.235 62.42 220.405 ;
     RECT  69.42 220.235 69.59 220.405 ;
     RECT  71.72 220.235 71.89 220.405 ;
     RECT  74.665 220.235 74.835 220.405 ;
     RECT  76.78 220.235 76.95 220.405 ;
     RECT  81.57 220.235 81.74 220.405 ;
     RECT  85.06 220.235 85.23 220.405 ;
     RECT  88.93 220.235 89.1 220.405 ;
     RECT  90.12 220.235 90.29 220.405 ;
     RECT  93.985 220.235 94.155 220.405 ;
     RECT  94.26 220.235 94.43 220.405 ;
     RECT  98.59 220.235 98.76 220.405 ;
     RECT  102.725 220.235 102.895 220.405 ;
     RECT  103.46 220.235 103.63 220.405 ;
     RECT  107.33 220.235 107.5 220.405 ;
     RECT  112.2 220.235 112.37 220.405 ;
     RECT  112.385 220.235 112.555 220.405 ;
     RECT  116.34 220.235 116.51 220.405 ;
     RECT  15.325 220.64 15.495 221.165 ;
     RECT  42.925 220.64 43.095 221.165 ;
     RECT  70.525 220.64 70.695 221.165 ;
     RECT  98.125 220.64 98.295 221.165 ;
     RECT  29.125 224.915 29.295 225.44 ;
     RECT  56.725 224.915 56.895 225.44 ;
     RECT  84.325 224.915 84.495 225.44 ;
     RECT  111.925 224.915 112.095 225.44 ;
     RECT  1.555 225.7 1.665 225.705 ;
     RECT  42.47 225.675 42.64 225.705 ;
     RECT  70.985 225.675 71.155 225.705 ;
     RECT  59.035 225.7 59.195 225.81 ;
     RECT  69.615 225.7 69.775 225.81 ;
     RECT  1.52 225.705 1.665 225.815 ;
     RECT  3.36 225.705 3.48 225.815 ;
     RECT  20.38 225.705 20.5 225.815 ;
     RECT  36.94 225.705 37.06 225.815 ;
     RECT  42.46 225.705 42.64 225.815 ;
     RECT  70.06 225.705 70.18 225.815 ;
     RECT  70.52 225.705 70.64 225.815 ;
     RECT  70.98 225.705 71.155 225.815 ;
     RECT  77.42 225.705 77.54 225.815 ;
     RECT  93.52 225.705 93.64 225.815 ;
     RECT  111.92 225.705 112.04 225.815 ;
     RECT  120.66 225.705 120.78 225.815 ;
     RECT  1.555 225.815 1.665 225.82 ;
     RECT  9.355 225.71 9.515 225.82 ;
     RECT  14.415 225.71 14.575 225.82 ;
     RECT  18.575 225.7 18.685 225.82 ;
     RECT  32.355 225.71 32.515 225.82 ;
     RECT  40.655 225.7 40.765 225.82 ;
     RECT  43.395 225.71 43.555 225.82 ;
     RECT  57.215 225.7 57.325 225.82 ;
     RECT  69.155 225.71 69.315 225.82 ;
     RECT  75.615 225.7 75.725 225.82 ;
     RECT  82.515 225.7 82.625 225.82 ;
     RECT  91.715 225.7 91.825 225.82 ;
     RECT  99.075 225.7 99.185 225.82 ;
     RECT  110.115 225.7 110.225 225.82 ;
     RECT  119.755 225.71 119.915 225.82 ;
     RECT  1.985 225.675 2.155 225.845 ;
     RECT  3.825 225.675 3.995 225.845 ;
     RECT  10.54 225.675 10.71 225.845 ;
     RECT  11.185 225.675 11.355 225.845 ;
     RECT  15.785 225.675 15.955 225.845 ;
     RECT  21.12 225.675 21.29 225.845 ;
     RECT  23.145 225.675 23.315 225.845 ;
     RECT  25.26 225.675 25.43 225.845 ;
     RECT  29.585 225.675 29.755 225.845 ;
     RECT  33.265 225.675 33.435 225.845 ;
     RECT  37.41 225.675 37.58 225.845 ;
     RECT  42.47 225.815 42.64 225.845 ;
     RECT  44.305 225.675 44.475 225.845 ;
     RECT  47.525 225.675 47.695 225.845 ;
     RECT  51.665 225.675 51.835 225.845 ;
     RECT  55.345 225.675 55.515 225.845 ;
     RECT  59.945 225.675 60.115 225.845 ;
     RECT  65.28 225.675 65.45 225.845 ;
     RECT  70.985 225.815 71.155 225.845 ;
     RECT  71.72 225.675 71.89 225.845 ;
     RECT  77.885 225.675 78.055 225.845 ;
     RECT  78.62 225.675 78.79 225.845 ;
     RECT  84.79 225.675 84.96 225.845 ;
     RECT  87.085 225.675 87.255 225.845 ;
     RECT  87.82 225.675 87.99 225.845 ;
     RECT  93.99 225.675 94.16 225.845 ;
     RECT  94.45 225.675 94.62 225.845 ;
     RECT  98.86 225.675 99.03 225.845 ;
     RECT  100.885 225.675 101.055 225.845 ;
     RECT  102.725 225.675 102.895 225.845 ;
     RECT  108.245 225.675 108.415 225.845 ;
     RECT  112.385 225.675 112.555 225.845 ;
     RECT  112.66 225.675 112.83 225.845 ;
     RECT  116.8 225.675 116.97 225.845 ;
     RECT  15.325 226.08 15.495 226.605 ;
     RECT  42.925 226.08 43.095 226.605 ;
     RECT  70.525 226.08 70.695 226.605 ;
     RECT  98.125 226.08 98.295 226.605 ;
     RECT  29.125 230.355 29.295 230.88 ;
     RECT  56.725 230.355 56.895 230.88 ;
     RECT  84.325 230.355 84.495 230.88 ;
     RECT  111.925 230.355 112.095 230.88 ;
     RECT  68.695 231.14 68.855 231.25 ;
     RECT  77.435 231.14 77.595 231.25 ;
     RECT  2.44 231.145 2.56 231.255 ;
     RECT  31.42 231.145 31.54 231.255 ;
     RECT  43.38 231.145 43.5 231.255 ;
     RECT  69.6 231.145 69.72 231.255 ;
     RECT  72.82 231.145 72.94 231.255 ;
     RECT  86.62 231.145 86.74 231.255 ;
     RECT  120.66 231.145 120.78 231.255 ;
     RECT  19.935 231.15 20.095 231.26 ;
     RECT  29.615 231.14 29.725 231.26 ;
     RECT  54.915 231.14 55.025 231.26 ;
     RECT  71.015 231.14 71.125 231.26 ;
     RECT  82.515 231.14 82.625 231.26 ;
     RECT  84.815 231.14 84.925 231.26 ;
     RECT  96.315 231.14 96.425 231.26 ;
     RECT  103.655 231.15 103.815 231.26 ;
     RECT  119.755 231.14 119.915 231.26 ;
     RECT  1.525 231.115 1.695 231.285 ;
     RECT  3.18 231.115 3.35 231.285 ;
     RECT  7.045 231.115 7.215 231.285 ;
     RECT  7.965 231.115 8.135 231.285 ;
     RECT  15.6 231.115 15.77 231.285 ;
     RECT  16.06 231.115 16.23 231.285 ;
     RECT  19.465 231.115 19.635 231.285 ;
     RECT  20.845 231.115 21.015 231.285 ;
     RECT  28.205 231.115 28.375 231.285 ;
     RECT  31.885 231.115 32.055 231.285 ;
     RECT  35.565 231.115 35.735 231.285 ;
     RECT  41.545 231.115 41.715 231.285 ;
     RECT  44.12 231.115 44.29 231.285 ;
     RECT  45.225 231.115 45.395 231.285 ;
     RECT  47.985 231.115 48.155 231.285 ;
     RECT  55.62 231.115 55.79 231.285 ;
     RECT  57.185 231.115 57.355 231.285 ;
     RECT  59.49 231.115 59.66 231.285 ;
     RECT  63.165 231.115 63.335 231.285 ;
     RECT  64.82 231.115 64.99 231.285 ;
     RECT  70.065 231.115 70.235 231.285 ;
     RECT  73.285 231.115 73.455 231.285 ;
     RECT  78.62 231.115 78.79 231.285 ;
     RECT  80.645 231.115 80.815 231.285 ;
     RECT  87.085 231.115 87.255 231.285 ;
     RECT  88.28 231.115 88.45 231.285 ;
     RECT  92.42 231.115 92.59 231.285 ;
     RECT  94.445 231.115 94.615 231.285 ;
     RECT  98.59 231.115 98.76 231.285 ;
     RECT  101.805 231.115 101.975 231.285 ;
     RECT  104.57 231.115 104.74 231.285 ;
     RECT  109.17 231.115 109.34 231.285 ;
     RECT  112.385 231.115 112.555 231.285 ;
     RECT  114.69 231.115 114.86 231.285 ;
     RECT  15.325 231.52 15.495 232.045 ;
     RECT  42.925 231.52 43.095 232.045 ;
     RECT  70.525 231.52 70.695 232.045 ;
     RECT  98.125 231.52 98.295 232.045 ;
     RECT  29.125 235.795 29.295 236.32 ;
     RECT  56.725 235.795 56.895 236.32 ;
     RECT  84.325 235.795 84.495 236.32 ;
     RECT  111.925 235.795 112.095 236.32 ;
     RECT  29.615 236.58 29.725 236.59 ;
     RECT  19.015 236.58 19.175 236.69 ;
     RECT  31.435 236.58 31.595 236.69 ;
     RECT  82.955 236.58 83.115 236.69 ;
     RECT  4.74 236.585 4.86 236.695 ;
     RECT  39.7 236.585 39.82 236.695 ;
     RECT  43.38 236.585 43.5 236.695 ;
     RECT  47.98 236.585 48.1 236.695 ;
     RECT  76.04 236.585 76.16 236.695 ;
     RECT  83.86 236.585 83.98 236.695 ;
     RECT  86.62 236.585 86.74 236.695 ;
     RECT  92.14 236.585 92.26 236.695 ;
     RECT  97.66 236.585 97.78 236.695 ;
     RECT  101.34 236.585 101.46 236.695 ;
     RECT  120.66 236.585 120.78 236.695 ;
     RECT  2.935 236.58 3.045 236.7 ;
     RECT  23.175 236.58 23.285 236.7 ;
     RECT  27.315 236.58 27.425 236.7 ;
     RECT  29.595 236.59 29.755 236.7 ;
     RECT  54.915 236.58 55.025 236.7 ;
     RECT  62.255 236.59 62.415 236.7 ;
     RECT  75.135 236.59 75.295 236.7 ;
     RECT  81.135 236.58 81.245 236.7 ;
     RECT  84.815 236.58 84.925 236.7 ;
     RECT  88.955 236.58 89.065 236.7 ;
     RECT  96.755 236.59 96.915 236.7 ;
     RECT  98.615 236.58 98.725 236.7 ;
     RECT  100.435 236.59 100.595 236.7 ;
     RECT  119.755 236.59 119.915 236.7 ;
     RECT  1.525 236.555 1.695 236.725 ;
     RECT  5.21 236.555 5.38 236.725 ;
     RECT  8.89 236.555 9.06 236.725 ;
     RECT  11.645 236.555 11.815 236.725 ;
     RECT  15.785 236.555 15.955 236.725 ;
     RECT  19.925 236.555 20.095 236.725 ;
     RECT  25.26 236.555 25.43 236.725 ;
     RECT  30.78 236.555 30.95 236.725 ;
     RECT  32.345 236.555 32.515 236.725 ;
     RECT  34.92 236.555 35.09 236.725 ;
     RECT  39.06 236.555 39.23 236.725 ;
     RECT  40.165 236.555 40.335 236.725 ;
     RECT  44.12 236.555 44.29 236.725 ;
     RECT  47.525 236.555 47.695 236.725 ;
     RECT  48.72 236.555 48.89 236.725 ;
     RECT  52.86 236.555 53.03 236.725 ;
     RECT  57.185 236.555 57.355 236.725 ;
     RECT  58.38 236.555 58.55 236.725 ;
     RECT  63.165 236.555 63.335 236.725 ;
     RECT  64.82 236.555 64.99 236.725 ;
     RECT  68.96 236.555 69.13 236.725 ;
     RECT  71.26 236.555 71.43 236.725 ;
     RECT  72.83 236.555 73 236.725 ;
     RECT  76.505 236.555 76.675 236.725 ;
     RECT  85.06 236.555 85.23 236.725 ;
     RECT  87.09 236.555 87.26 236.725 ;
     RECT  90.77 236.555 90.94 236.725 ;
     RECT  92.88 236.555 93.05 236.725 ;
     RECT  100.885 236.555 101.055 236.725 ;
     RECT  101.81 236.555 101.98 236.725 ;
     RECT  108.245 236.555 108.415 236.725 ;
     RECT  112.385 236.555 112.555 236.725 ;
     RECT  113.305 236.555 113.475 236.725 ;
     RECT  15.325 236.96 15.495 237.485 ;
     RECT  29.125 236.96 29.295 237.485 ;
     RECT  42.925 236.96 43.095 237.485 ;
     RECT  56.725 236.96 56.895 237.485 ;
     RECT  70.525 236.96 70.695 237.485 ;
     RECT  84.325 236.96 84.495 237.485 ;
     RECT  98.125 236.96 98.295 237.485 ;
     RECT  111.925 236.96 112.095 237.485 ;
    LAYER li1 ;
     RECT  1.38 2.635 120.98 239.445 ;
    LAYER met1 ;
     RECT  -6.62 5.2 1.08 239.6 ;
     RECT  1.08 2.14 6.14 239.6 ;
     RECT  6.14 2.14 13.96 240.62 ;
     RECT  13.96 2.14 18.7 240.96 ;
     RECT  18.7 2.48 73.9 240.96 ;
     RECT  73.9 2.48 78.96 240.28 ;
     RECT  78.96 2.48 85.72 239.6 ;
     RECT  85.72 0.78 109.78 239.6 ;
     RECT  109.78 1.46 120.36 239.6 ;
     RECT  120.36 2.48 124.98 239.6 ;
     RECT  124.98 5.2 128.98 239.6 ;
    LAYER met2 ;
     RECT  85.72 0.78 85.86 1.46 ;
     RECT  109.64 0.78 109.78 1.46 ;
     RECT  85.72 1.46 94.14 1.8 ;
     RECT  105.04 1.46 120.36 2.535 ;
     RECT  18.56 2.14 18.7 3.5 ;
     RECT  85.72 1.8 95.52 3.5 ;
     RECT  18.56 3.5 27.44 3.84 ;
     RECT  38.8 3.5 38.94 3.84 ;
     RECT  56.74 3.5 56.88 3.84 ;
     RECT  76.06 3.5 95.52 3.84 ;
     RECT  6.6 3.84 6.74 4.18 ;
     RECT  18.56 3.84 43.54 4.18 ;
     RECT  54.44 3.84 95.52 4.18 ;
     RECT  105.04 2.535 124.92 4.18 ;
     RECT  54.44 4.18 124.92 4.86 ;
     RECT  1.54 4.18 43.54 5.255 ;
     RECT  53.06 4.86 124.92 5.255 ;
     RECT  -6.56 5.255 43.54 6.22 ;
     RECT  53.06 5.255 128.92 6.22 ;
     RECT  -6.56 6.22 128.92 236.825 ;
     RECT  -6.56 236.825 117.6 237.22 ;
     RECT  -6.56 237.22 80.34 237.56 ;
     RECT  90.32 237.22 117.6 237.56 ;
     RECT  90.32 237.56 112.54 237.9 ;
     RECT  -6.56 237.56 78.96 238.24 ;
     RECT  56.74 238.24 58.26 238.58 ;
     RECT  93.08 237.9 110.7 238.58 ;
     RECT  -6.56 238.24 38.02 238.92 ;
     RECT  104.58 238.58 110.7 238.92 ;
     RECT  -6.56 238.92 26.52 239.545 ;
     RECT  127.04 236.825 128.92 239.545 ;
     RECT  2.92 239.545 26.52 240.28 ;
     RECT  68.7 238.24 78.96 240.28 ;
     RECT  2.92 240.28 20.08 240.62 ;
     RECT  68.7 240.28 73.9 240.62 ;
     RECT  13.96 240.62 20.08 240.96 ;
     RECT  73.76 240.62 73.9 240.96 ;
     RECT  2.92 240.62 3.98 242.19 ;
     RECT  93.08 238.58 93.22 242.19 ;
     RECT  106.88 238.92 110.7 242.19 ;
    LAYER met3 ;
     RECT  -6.62 -5.28 -6.61 -3.28 ;
     RECT  -6.62 245.36 -6.61 247.36 ;
     RECT  -6.61 -5.28 -4.63 247.36 ;
     RECT  -4.63 108.99 6.13 145.33 ;
     RECT  -4.63 -5.28 9.74 17.49 ;
     RECT  -4.63 83.83 9.74 84.13 ;
     RECT  9.74 72.27 11.8 84.13 ;
     RECT  6.13 108.99 11.8 129.69 ;
     RECT  -4.63 192.63 12.5 214.01 ;
     RECT  -4.63 230.03 12.5 247.36 ;
     RECT  11.12 175.63 12.96 175.93 ;
     RECT  6.13 143.67 13.95 145.33 ;
     RECT  11.8 72.27 20.32 129.69 ;
     RECT  13.95 143.67 20.32 143.97 ;
     RECT  12.96 175.63 20.32 178.65 ;
     RECT  12.5 192.63 20.32 247.36 ;
     RECT  20.32 72.27 20.62 143.97 ;
     RECT  20.32 175.63 20.85 247.36 ;
     RECT  9.74 -5.28 26.14 20.21 ;
     RECT  20.62 72.27 27.22 143.29 ;
     RECT  26.14 17.19 28.14 20.21 ;
     RECT  20.85 175.63 28.14 226.25 ;
     RECT  28.14 17.19 28.83 25.65 ;
     RECT  28.83 17.19 29.06 30.41 ;
     RECT  27.22 58.67 32.12 143.29 ;
     RECT  32.12 61.39 34.58 143.29 ;
     RECT  28.14 165.43 34.58 226.25 ;
     RECT  29.06 17.19 39.94 34.49 ;
     RECT  34.58 61.39 41.32 226.25 ;
     RECT  41.32 61.39 41.78 72.57 ;
     RECT  41.32 87.91 41.94 226.25 ;
     RECT  20.85 241.36 41.94 247.36 ;
     RECT  41.94 87.91 42.7 247.36 ;
     RECT  42.7 87.91 43.62 137.85 ;
     RECT  43.62 87.91 45.46 96.37 ;
     RECT  45.46 87.91 45.92 88.21 ;
     RECT  39.94 17.19 46.38 18.17 ;
     RECT  42.7 156.59 46.84 247.36 ;
     RECT  41.78 61.39 47.68 61.69 ;
     RECT  39.94 34.19 47.7 34.49 ;
     RECT  47.7 34.19 48.45 35.17 ;
     RECT  47.68 55.27 48.45 61.69 ;
     RECT  48.45 34.87 48.68 35.17 ;
     RECT  43.62 110.35 49.14 137.85 ;
     RECT  46.84 157.95 55.12 247.36 ;
     RECT  55.28 81.11 56.66 81.41 ;
     RECT  56.66 79.07 60.8 81.41 ;
     RECT  48.45 61.39 62.87 61.69 ;
     RECT  62.87 61.39 63.17 62.37 ;
     RECT  46.38 17.19 67.08 17.49 ;
     RECT  63.17 62.07 67.7 62.37 ;
     RECT  67.7 62.07 71.38 63.73 ;
     RECT  60.8 79.07 71.38 90.25 ;
     RECT  49.14 111.03 71.38 137.85 ;
     RECT  60.8 151.83 71.38 152.13 ;
     RECT  71.38 62.07 75.75 90.25 ;
     RECT  71.38 111.03 75.75 152.13 ;
     RECT  75.75 62.07 82.49 152.13 ;
     RECT  75.52 41.67 83.34 41.97 ;
     RECT  82.49 62.07 83.64 97.05 ;
     RECT  55.12 172.23 86.79 247.36 ;
     RECT  82.49 111.03 87.09 152.13 ;
     RECT  81.96 19.91 89.31 20.21 ;
     RECT  87.09 117.15 89.32 152.13 ;
     RECT  86.79 166.79 89.32 247.36 ;
     RECT  89.31 19.23 89.55 20.21 ;
     RECT  89.55 19.23 91.16 20.89 ;
     RECT  83.34 34.87 92.61 41.97 ;
     RECT  92.61 34.87 93.08 40.61 ;
     RECT  91.16 17.87 96.98 20.89 ;
     RECT  89.32 117.15 97.44 247.36 ;
     RECT  83.64 67.51 98.06 97.05 ;
     RECT  98.06 58.67 100.82 97.05 ;
     RECT  97.44 117.15 100.82 117.45 ;
     RECT  96.98 17.87 101.74 18.17 ;
     RECT  97.44 131.43 103.42 247.36 ;
     RECT  103.42 131.43 103.65 214.69 ;
     RECT  100.82 58.67 104.04 117.45 ;
     RECT  103.42 232.75 105.26 247.36 ;
     RECT  26.14 -5.28 105.42 0.72 ;
     RECT  101.74 15.15 105.42 18.17 ;
     RECT  103.65 131.43 105.72 210.61 ;
     RECT  93.08 34.87 107.26 35.17 ;
     RECT  105.72 175.63 108.02 210.61 ;
     RECT  104.04 57.31 108.48 117.45 ;
     RECT  108.02 180.39 108.94 210.61 ;
     RECT  105.42 -5.28 112.78 18.17 ;
     RECT  107.26 33.51 112.78 35.17 ;
     RECT  112.78 -5.28 122.99 35.17 ;
     RECT  108.48 58.67 122.99 117.45 ;
     RECT  105.72 131.43 122.99 158.25 ;
     RECT  108.94 180.39 122.99 209.93 ;
     RECT  105.26 241.36 122.99 247.36 ;
     RECT  122.99 -5.28 128.97 247.36 ;
     RECT  128.97 -5.28 128.98 -3.28 ;
     RECT  128.97 245.36 128.98 247.36 ;
    LAYER met4 ;
     RECT  -6.62 -5.28 -4.62 -1.28 ;
     RECT  126.98 -5.28 128.98 -1.28 ;
     RECT  28.83 19.91 29.13 30.41 ;
     RECT  89.55 19.23 89.85 40.31 ;
     RECT  48.15 34.87 48.45 55.57 ;
     RECT  89.55 40.31 92.61 67.51 ;
     RECT  -6.62 -1.28 -0.62 72.27 ;
     RECT  65.63 62.07 65.93 75.67 ;
     RECT  89.55 67.51 94.45 75.67 ;
     RECT  65.63 75.67 95.37 95.39 ;
     RECT  -6.62 72.27 12.57 97.05 ;
     RECT  65.63 95.39 97.21 110.35 ;
     RECT  47.23 110.35 97.21 123.95 ;
     RECT  41.71 123.95 97.21 144.35 ;
     RECT  40.79 144.35 97.21 145.03 ;
     RECT  40.79 145.03 98.13 151.83 ;
     RECT  35.27 151.83 103.65 186.81 ;
     RECT  35.27 186.81 75.13 193.31 ;
     RECT  20.55 193.31 75.13 193.61 ;
     RECT  20.55 193.61 42.93 209.93 ;
     RECT  74.83 193.61 75.13 214.01 ;
     RECT  95.07 186.81 103.65 214.69 ;
     RECT  95.07 214.69 95.37 221.49 ;
     RECT  20.55 209.93 35.57 225.57 ;
     RECT  20.55 225.57 20.85 233.05 ;
     RECT  -6.62 97.05 -0.62 243.36 ;
     RECT  122.98 -1.28 128.98 243.36 ;
     RECT  -6.62 243.36 -4.62 247.36 ;
     RECT  126.98 243.36 128.98 247.36 ;
  END
END fifo
END LIBRARY
