VERSION 5.7 ;
NAMESCASESENSITIVE ON ;
BUSBITCHARS "[]" ;
DIVIDERCHAR "/" ;

PROPERTYDEFINITIONS
    LAYER LEF58_TYPE STRING ;
END PROPERTYDEFINITIONS

UNITS
    DATABASE MICRONS 1000 ;
END UNITS
USEMINSPACING OBS OFF ;
MANUFACTURINGGRID 0.005 ;

LAYER nwell
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE NWELL ;" ;
END nwell

LAYER pwell
    TYPE MASTERSLICE ;
    PROPERTY LEF58_TYPE "TYPE PWELL ;" ;
END pwell

LAYER li1
    TYPE ROUTING ;
    PITCH 0.46 ;
    WIDTH 0.17 ;
    AREA 0.0561 ;
    THICKNESS 0.1 ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 0.170 ;
    ANTENNADIFFSIDEAREARATIO  PWL ( ( 0 75 ) ( 0.0125 75 ) ( 0.0225 85.125 ) ( 22.5 10200 ) ) ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 12.199200031 ;
    CAPACITANCE CPERSQDIST 0.00088176470459 ;
END li1

LAYER mcon
    TYPE CUT ;
    WIDTH 0.17 ;
    SPACING 0.19  ;
    ANTENNADIFFAREARATIO  PWL ( ( 0 3 ) ( 0.0125 3 ) ( 0.0225 3.405 ) ( 22.5 408 ) ) ;
    RESISTANCE 9.249146 ;
END mcon

LAYER met1
    TYPE ROUTING ;
    PITCH 0.34 ;
    WIDTH 0.14 ;
    AREA 0.083 ;
    THICKNESS 0.35 ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 0.140
  WIDTH 3.000	 0.280 ;
    MINENCLOSEDAREA 0.14 ;
    ANTENNADIFFSIDEAREARATIO  PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.12500600032 ;
    CAPACITANCE CPERSQDIST 0.0012312499982 ;
END met1

LAYER via
    TYPE CUT ;
    WIDTH 0.15 ;
    SPACING 0.17  ;
    ANTENNADIFFAREARATIO  PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
    RESISTANCE 4.5 ;
END via

LAYER met2
    TYPE ROUTING ;
    PITCH 0.46 ;
    WIDTH 0.14 ;
    AREA 0.0676 ;
    THICKNESS 0.35 ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 0.140
  WIDTH 3.000	 0.280 ;
    MINENCLOSEDAREA 0.14 ;
    ANTENNADIFFSIDEAREARATIO  PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.12500600032 ;
    CAPACITANCE CPERSQDIST 0.00097309285571 ;
END met2

LAYER via2
    TYPE CUT ;
    WIDTH 0.2 ;
    SPACING 0.2  ;
    ANTENNADIFFAREARATIO  PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
    RESISTANCE 3.368786 ;
END via2

LAYER met3
    TYPE ROUTING ;
    PITCH 0.68 ;
    WIDTH 0.3 ;
    AREA 0.24 ;
    THICKNESS 0.8 ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 0.300
  WIDTH 3.000	 0.400 ;
    ANTENNADIFFSIDEAREARATIO  PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.047010000119 ;
    CAPACITANCE CPERSQDIST 0.00071653999895 ;
END met3

LAYER via3
    TYPE CUT ;
    WIDTH 0.2 ;
    SPACING 0.2  ;
    ANTENNADIFFAREARATIO  PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
    RESISTANCE 0.376635 ;
END via3

LAYER met4
    TYPE ROUTING ;
    PITCH 0.92 ;
    WIDTH 0.3 ;
    AREA 0.24 ;
    THICKNESS 0.8 ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 0.300
  WIDTH 3.000	 0.400 ;
    ANTENNADIFFSIDEAREARATIO  PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
    DIRECTION VERTICAL ;
    RESISTANCE RPERSQ 0.047010000119 ;
    CAPACITANCE CPERSQDIST 0.00049375999927 ;
END met4

LAYER via4
    TYPE CUT ;
    WIDTH 0.8 ;
    SPACING 0.8  ;
    ANTENNADIFFAREARATIO  PWL ( ( 0 6 ) ( 0.0125 6 ) ( 0.0225 6.81 ) ( 22.5 816 ) ) ;
    RESISTANCE 0.0058 ;
END via4

LAYER met5
    TYPE ROUTING ;
    PITCH 3.4 ;
    WIDTH 1.6 ;
    AREA 4 ;
    THICKNESS 1.2 ;
SPACINGTABLE
  PARALLELRUNLENGTH 0.000
  WIDTH 0.000	 1.600 ;
    ANTENNADIFFSIDEAREARATIO  PWL ( ( 0 400 ) ( 0.0125 400 ) ( 0.0225 2609 ) ( 22.5 11600 ) ) ;
    DIRECTION HORIZONTAL ;
    RESISTANCE RPERSQ 0.028496000072 ;
    CAPACITANCE CPERSQDIST 9.6304374858e-05 ;
END met5

VIA L1M1_PR DEFAULT
    LAYER mcon ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER li1 ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER met1 ;
      RECT  -0.145 -0.115 0.145 0.115 ;
END L1M1_PR

VIA L1M1_PR_R DEFAULT
    LAYER mcon ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER li1 ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER met1 ;
      RECT  -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_R

VIA L1M1_PR_M DEFAULT
    LAYER mcon ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER li1 ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER met1 ;
      RECT  -0.115 -0.145 0.115 0.145 ;
END L1M1_PR_M

VIA L1M1_PR_MR DEFAULT
    LAYER mcon ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER li1 ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER met1 ;
      RECT  -0.145 -0.115 0.145 0.115 ;
END L1M1_PR_MR

VIA L1M1_PR_C DEFAULT
    LAYER mcon ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER li1 ;
      RECT  -0.085 -0.085 0.085 0.085 ;
    LAYER met1 ;
      RECT  -0.145 -0.145 0.145 0.145 ;
END L1M1_PR_C

VIA M1M2_PR DEFAULT
    LAYER via ;
      RECT  -0.075 -0.075 0.075 0.075 ;
    LAYER met1 ;
      RECT  -0.16 -0.13 0.16 0.13 ;
    LAYER met2 ;
      RECT  -0.13 -0.16 0.13 0.16 ;
END M1M2_PR

VIA M1M2_PR_R DEFAULT
    LAYER via ;
      RECT  -0.075 -0.075 0.075 0.075 ;
    LAYER met1 ;
      RECT  -0.13 -0.16 0.13 0.16 ;
    LAYER met2 ;
      RECT  -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_R

VIA M1M2_PR_M DEFAULT
    LAYER via ;
      RECT  -0.075 -0.075 0.075 0.075 ;
    LAYER met1 ;
      RECT  -0.16 -0.13 0.16 0.13 ;
    LAYER met2 ;
      RECT  -0.16 -0.13 0.16 0.13 ;
END M1M2_PR_M

VIA M1M2_PR_MR DEFAULT
    LAYER via ;
      RECT  -0.075 -0.075 0.075 0.075 ;
    LAYER met1 ;
      RECT  -0.13 -0.16 0.13 0.16 ;
    LAYER met2 ;
      RECT  -0.13 -0.16 0.13 0.16 ;
END M1M2_PR_MR

VIA M1M2_PR_C DEFAULT
    LAYER via ;
      RECT  -0.075 -0.075 0.075 0.075 ;
    LAYER met1 ;
      RECT  -0.16 -0.16 0.16 0.16 ;
    LAYER met2 ;
      RECT  -0.16 -0.16 0.16 0.16 ;
END M1M2_PR_C

VIA M2M3_PR DEFAULT
    LAYER via2 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met2 ;
      RECT  -0.14 -0.185 0.14 0.185 ;
    LAYER met3 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M2M3_PR

VIA M2M3_PR_R DEFAULT
    LAYER via2 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met2 ;
      RECT  -0.185 -0.14 0.185 0.14 ;
    LAYER met3 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_R

VIA M2M3_PR_M DEFAULT
    LAYER via2 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met2 ;
      RECT  -0.14 -0.185 0.14 0.185 ;
    LAYER met3 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_M

VIA M2M3_PR_MR DEFAULT
    LAYER via2 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met2 ;
      RECT  -0.185 -0.14 0.185 0.14 ;
    LAYER met3 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_MR

VIA M2M3_PR_C DEFAULT
    LAYER via2 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met2 ;
      RECT  -0.185 -0.185 0.185 0.185 ;
    LAYER met3 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M2M3_PR_C

VIA M3M4_PR DEFAULT
    LAYER via3 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met3 ;
      RECT  -0.19 -0.16 0.19 0.16 ;
    LAYER met4 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M3M4_PR

VIA M3M4_PR_R DEFAULT
    LAYER via3 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met3 ;
      RECT  -0.16 -0.19 0.16 0.19 ;
    LAYER met4 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_R

VIA M3M4_PR_M DEFAULT
    LAYER via3 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met3 ;
      RECT  -0.19 -0.16 0.19 0.16 ;
    LAYER met4 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_M

VIA M3M4_PR_MR DEFAULT
    LAYER via3 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met3 ;
      RECT  -0.16 -0.19 0.16 0.19 ;
    LAYER met4 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_MR

VIA M3M4_PR_C DEFAULT
    LAYER via3 ;
      RECT  -0.1 -0.1 0.1 0.1 ;
    LAYER met3 ;
      RECT  -0.19 -0.19 0.19 0.19 ;
    LAYER met4 ;
      RECT  -0.165 -0.165 0.165 0.165 ;
END M3M4_PR_C

VIA M4M5_PR DEFAULT
    LAYER via4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
    LAYER met4 ;
      RECT  -0.59 -0.59 0.59 0.59 ;
    LAYER met5 ;
      RECT  -0.71 -0.71 0.71 0.71 ;
END M4M5_PR

VIA M4M5_PR_R DEFAULT
    LAYER via4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
    LAYER met4 ;
      RECT  -0.59 -0.59 0.59 0.59 ;
    LAYER met5 ;
      RECT  -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_R

VIA M4M5_PR_M DEFAULT
    LAYER via4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
    LAYER met4 ;
      RECT  -0.59 -0.59 0.59 0.59 ;
    LAYER met5 ;
      RECT  -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_M

VIA M4M5_PR_MR DEFAULT
    LAYER via4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
    LAYER met4 ;
      RECT  -0.59 -0.59 0.59 0.59 ;
    LAYER met5 ;
      RECT  -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_MR

VIA M4M5_PR_C DEFAULT
    LAYER via4 ;
      RECT  -0.4 -0.4 0.4 0.4 ;
    LAYER met4 ;
      RECT  -0.59 -0.59 0.59 0.59 ;
    LAYER met5 ;
      RECT  -0.71 -0.71 0.71 0.71 ;
END M4M5_PR_C

VIARULE L1M1_PR GENERATE 
    LAYER li1 ;
      ENCLOSURE 0 0 ;
    LAYER met1 ;
      ENCLOSURE 0.06 0.03 ;
    LAYER mcon ;
      RECT  -0.085 -0.085  0.085 0.085  ;
      SPACING 0.36 BY 0.36 ;
END L1M1_PR

VIARULE L1M1_PR_R GENERATE 
    LAYER li1 ;
      ENCLOSURE 0 0 ;
    LAYER met1 ;
      ENCLOSURE 0.03 0.06 ;
    LAYER mcon ;
      RECT  -0.085 -0.085  0.085 0.085  ;
      SPACING 0.36 BY 0.36 ;
END L1M1_PR_R

VIARULE L1M1_PR_M GENERATE 
    LAYER li1 ;
      ENCLOSURE 0 0 ;
    LAYER met1 ;
      ENCLOSURE 0.03 0.06 ;
    LAYER mcon ;
      RECT  -0.085 -0.085  0.085 0.085  ;
      SPACING 0.36 BY 0.36 ;
END L1M1_PR_M

VIARULE L1M1_PR_MR GENERATE 
    LAYER li1 ;
      ENCLOSURE 0 0 ;
    LAYER met1 ;
      ENCLOSURE 0.06 0.03 ;
    LAYER mcon ;
      RECT  -0.085 -0.085  0.085 0.085  ;
      SPACING 0.36 BY 0.36 ;
END L1M1_PR_MR

VIARULE L1M1_PR_C GENERATE 
    LAYER li1 ;
      ENCLOSURE 0 0 ;
    LAYER met1 ;
      ENCLOSURE 0.06 0.06 ;
    LAYER mcon ;
      RECT  -0.085 -0.085  0.085 0.085  ;
      SPACING 0.36 BY 0.36 ;
END L1M1_PR_C

VIARULE M1M2_PR GENERATE 
    LAYER met1 ;
      ENCLOSURE 0.085 0.055 ;
    LAYER met2 ;
      ENCLOSURE 0.055 0.085 ;
    LAYER via ;
      RECT  -0.075 -0.075  0.075 0.075  ;
      SPACING 0.32 BY 0.32 ;
END M1M2_PR

VIARULE M1M2_PR_R GENERATE 
    LAYER met1 ;
      ENCLOSURE 0.055 0.085 ;
    LAYER met2 ;
      ENCLOSURE 0.085 0.055 ;
    LAYER via ;
      RECT  -0.075 -0.075  0.075 0.075  ;
      SPACING 0.32 BY 0.32 ;
END M1M2_PR_R

VIARULE M1M2_PR_M GENERATE 
    LAYER met1 ;
      ENCLOSURE 0.085 0.055 ;
    LAYER met2 ;
      ENCLOSURE 0.085 0.055 ;
    LAYER via ;
      RECT  -0.075 -0.075  0.075 0.075  ;
      SPACING 0.32 BY 0.32 ;
END M1M2_PR_M

VIARULE M1M2_PR_MR GENERATE 
    LAYER met1 ;
      ENCLOSURE 0.055 0.085 ;
    LAYER met2 ;
      ENCLOSURE 0.055 0.085 ;
    LAYER via ;
      RECT  -0.075 -0.075  0.075 0.075  ;
      SPACING 0.32 BY 0.32 ;
END M1M2_PR_MR

VIARULE M1M2_PR_C GENERATE 
    LAYER met1 ;
      ENCLOSURE 0.085 0.085 ;
    LAYER met2 ;
      ENCLOSURE 0.085 0.085 ;
    LAYER via ;
      RECT  -0.075 -0.075  0.075 0.075  ;
      SPACING 0.32 BY 0.32 ;
END M1M2_PR_C

VIARULE M2M3_PR GENERATE 
    LAYER met2 ;
      ENCLOSURE 0.04 0.085 ;
    LAYER met3 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via2 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M2M3_PR

VIARULE M2M3_PR_R GENERATE 
    LAYER met2 ;
      ENCLOSURE 0.085 0.04 ;
    LAYER met3 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via2 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M2M3_PR_R

VIARULE M2M3_PR_M GENERATE 
    LAYER met2 ;
      ENCLOSURE 0.04 0.085 ;
    LAYER met3 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via2 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M2M3_PR_M

VIARULE M2M3_PR_MR GENERATE 
    LAYER met2 ;
      ENCLOSURE 0.085 0.04 ;
    LAYER met3 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via2 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M2M3_PR_MR

VIARULE M2M3_PR_C GENERATE 
    LAYER met2 ;
      ENCLOSURE 0.085 0.085 ;
    LAYER met3 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via2 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M2M3_PR_C

VIARULE M3M4_PR GENERATE 
    LAYER met3 ;
      ENCLOSURE 0.09 0.06 ;
    LAYER met4 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via3 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M3M4_PR

VIARULE M3M4_PR_R GENERATE 
    LAYER met3 ;
      ENCLOSURE 0.06 0.09 ;
    LAYER met4 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via3 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M3M4_PR_R

VIARULE M3M4_PR_M GENERATE 
    LAYER met3 ;
      ENCLOSURE 0.09 0.06 ;
    LAYER met4 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via3 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M3M4_PR_M

VIARULE M3M4_PR_MR GENERATE 
    LAYER met3 ;
      ENCLOSURE 0.06 0.09 ;
    LAYER met4 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via3 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M3M4_PR_MR

VIARULE M3M4_PR_C GENERATE 
    LAYER met3 ;
      ENCLOSURE 0.09 0.09 ;
    LAYER met4 ;
      ENCLOSURE 0.065 0.065 ;
    LAYER via3 ;
      RECT  -0.1 -0.1  0.1 0.1  ;
      SPACING 0.4 BY 0.4 ;
END M3M4_PR_C

VIARULE M4M5_PR GENERATE 
    LAYER met4 ;
      ENCLOSURE 0.19 0.19 ;
    LAYER met5 ;
      ENCLOSURE 0.31 0.31 ;
    LAYER via4 ;
      RECT  -0.4 -0.4  0.4 0.4  ;
      SPACING 1.6 BY 1.6 ;
END M4M5_PR

VIARULE M4M5_PR_R GENERATE 
    LAYER met4 ;
      ENCLOSURE 0.19 0.19 ;
    LAYER met5 ;
      ENCLOSURE 0.31 0.31 ;
    LAYER via4 ;
      RECT  -0.4 -0.4  0.4 0.4  ;
      SPACING 1.6 BY 1.6 ;
END M4M5_PR_R

VIARULE M4M5_PR_M GENERATE 
    LAYER met4 ;
      ENCLOSURE 0.19 0.19 ;
    LAYER met5 ;
      ENCLOSURE 0.31 0.31 ;
    LAYER via4 ;
      RECT  -0.4 -0.4  0.4 0.4  ;
      SPACING 1.6 BY 1.6 ;
END M4M5_PR_M

VIARULE M4M5_PR_MR GENERATE 
    LAYER met4 ;
      ENCLOSURE 0.19 0.19 ;
    LAYER met5 ;
      ENCLOSURE 0.31 0.31 ;
    LAYER via4 ;
      RECT  -0.4 -0.4  0.4 0.4  ;
      SPACING 1.6 BY 1.6 ;
END M4M5_PR_MR

VIARULE M4M5_PR_C GENERATE 
    LAYER met4 ;
      ENCLOSURE 0.19 0.19 ;
    LAYER met5 ;
      ENCLOSURE 0.31 0.31 ;
    LAYER via4 ;
      RECT  -0.4 -0.4  0.4 0.4  ;
      SPACING 1.6 BY 1.6 ;
END M4M5_PR_C
SITE unithd
    CLASS CORE ;
    SYMMETRY Y ;
    SIZE 0.46 BY 2.72 ;
END unithd
SITE unithddbl
    CLASS CORE ;
    SYMMETRY Y ;
    SIZE 0.46 BY 5.44 ;
END unithddbl
END LIBRARY
